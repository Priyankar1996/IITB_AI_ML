-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_50_load_0_ack_1 : boolean;
  signal ptr_deref_38_load_0_req_0 : boolean;
  signal ptr_deref_38_load_0_ack_0 : boolean;
  signal ptr_deref_38_load_0_req_1 : boolean;
  signal ptr_deref_38_load_0_ack_1 : boolean;
  signal ptr_deref_50_load_0_req_0 : boolean;
  signal ptr_deref_50_load_0_ack_0 : boolean;
  signal ptr_deref_50_load_0_req_1 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal ptr_deref_62_load_0_req_0 : boolean;
  signal ptr_deref_62_load_0_ack_0 : boolean;
  signal ptr_deref_62_load_0_req_1 : boolean;
  signal ptr_deref_62_load_0_ack_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal if_stmt_91_branch_req_0 : boolean;
  signal if_stmt_91_branch_ack_1 : boolean;
  signal if_stmt_91_branch_ack_0 : boolean;
  signal type_cast_110_inst_req_0 : boolean;
  signal type_cast_110_inst_ack_0 : boolean;
  signal type_cast_110_inst_req_1 : boolean;
  signal type_cast_110_inst_ack_1 : boolean;
  signal array_obj_ref_145_index_offset_req_0 : boolean;
  signal array_obj_ref_145_index_offset_ack_0 : boolean;
  signal array_obj_ref_145_index_offset_req_1 : boolean;
  signal array_obj_ref_145_index_offset_ack_1 : boolean;
  signal addr_of_146_final_reg_req_0 : boolean;
  signal addr_of_146_final_reg_ack_0 : boolean;
  signal addr_of_146_final_reg_req_1 : boolean;
  signal addr_of_146_final_reg_ack_1 : boolean;
  signal ptr_deref_150_load_0_req_0 : boolean;
  signal ptr_deref_150_load_0_ack_0 : boolean;
  signal ptr_deref_150_load_0_req_1 : boolean;
  signal ptr_deref_150_load_0_ack_1 : boolean;
  signal type_cast_154_inst_req_0 : boolean;
  signal type_cast_154_inst_ack_0 : boolean;
  signal type_cast_154_inst_req_1 : boolean;
  signal type_cast_154_inst_ack_1 : boolean;
  signal type_cast_174_inst_req_0 : boolean;
  signal type_cast_174_inst_ack_0 : boolean;
  signal type_cast_174_inst_req_1 : boolean;
  signal type_cast_174_inst_ack_1 : boolean;
  signal type_cast_184_inst_req_0 : boolean;
  signal type_cast_184_inst_ack_0 : boolean;
  signal type_cast_184_inst_req_1 : boolean;
  signal type_cast_184_inst_ack_1 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal type_cast_204_inst_req_0 : boolean;
  signal type_cast_204_inst_ack_0 : boolean;
  signal type_cast_204_inst_req_1 : boolean;
  signal type_cast_204_inst_ack_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal type_cast_224_inst_req_0 : boolean;
  signal type_cast_224_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_226_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_229_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_232_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_235_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_238_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_241_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_244_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_247_inst_ack_1 : boolean;
  signal if_stmt_261_branch_req_0 : boolean;
  signal if_stmt_261_branch_ack_1 : boolean;
  signal if_stmt_261_branch_ack_0 : boolean;
  signal phi_stmt_133_req_0 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal phi_stmt_133_req_1 : boolean;
  signal phi_stmt_133_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(68);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (86) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_27/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/branch_block_stmt_27__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/cr
      -- 
    rr_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_38_load_0_req_0); -- 
    cr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_38_load_0_req_1); -- 
    rr_139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_50_load_0_req_0); -- 
    cr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_50_load_0_req_1); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_62_load_0_req_0); -- 
    cr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => ptr_deref_62_load_0_req_1); -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => type_cast_76_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Sample/word_access_start/word_0/ra
      -- 
    ra_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_38_load_0_ack_0, ack => sendOutput_CP_26_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_38_Update/ptr_deref_38_Merge/merge_ack
      -- 
    ca_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_38_load_0_ack_1, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Sample/word_access_start/word_0/ra
      -- 
    ra_140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_50_load_0_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/ptr_deref_50_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_50_Update/word_access_complete/word_0/$exit
      -- 
    ca_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_50_load_0_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Sample/word_access_start/word_0/ra
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_62_load_0_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/ptr_deref_62_Update/ptr_deref_62_Merge/merge_ack
      -- 
    ca_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_62_load_0_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/rr
      -- 
    rr_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(7), ack => type_cast_76_inst_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(6) & sendOutput_CP_26_elements(4) & sendOutput_CP_26_elements(2);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Sample/ra
      -- 
    ra_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => sendOutput_CP_26_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (13) 
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90__exit__
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91__entry__
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/$exit
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_27/assign_stmt_35_to_assign_stmt_90/type_cast_76_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_27/R_cmp77_92_place
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/if_stmt_91_else_link/$entry
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => sendOutput_CP_26_elements(9)); -- 
    branch_req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(9), ack => if_stmt_91_branch_req_0); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	68 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_27/if_stmt_91_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_27/if_stmt_91_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_27/entry_forx_xend
      -- CP-element group 10: 	 branch_block_stmt_27/entry_forx_xend_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_27/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_91_branch_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (18) 
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97__exit__
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130__entry__
      -- CP-element group 11: 	 branch_block_stmt_27/if_stmt_91_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_27/if_stmt_91_else_link/else_choice_transition
      -- CP-element group 11: 	 branch_block_stmt_27/entry_bbx_xnph
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_update_start_
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_27/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_27/merge_stmt_97_PhiAck/dummy
      -- 
    else_choice_transition_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_91_branch_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_110_inst_req_0); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(11), ack => type_cast_110_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_0, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  place  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	62 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130__exit__
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/$exit
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_27/assign_stmt_102_to_assign_stmt_130/type_cast_110_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/$entry
      -- CP-element group 13: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$entry
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_1, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	59 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_sample_complete
      -- CP-element group 14: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/ack
      -- 
    ack_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_145_index_offset_ack_0, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	67 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (11) 
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/ack
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/$entry
      -- CP-element group 15: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/req
      -- 
    ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_145_index_offset_ack_1, ack => sendOutput_CP_26_elements(15)); -- 
    req_299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(15), ack => addr_of_146_final_reg_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/$exit
      -- CP-element group 16: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_request/ack
      -- 
    ack_300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_146_final_reg_ack_0, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (24) 
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_address_resized
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/base_resize_req
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_addr_resize/base_resize_ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/$exit
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/root_register_req
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_word_addrgen/root_register_ack
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/$entry
      -- CP-element group 17: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/rr
      -- 
    ack_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_146_final_reg_ack_1, ack => sendOutput_CP_26_elements(17)); -- 
    rr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(17), ack => ptr_deref_150_load_0_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/$exit
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Sample/word_access_start/word_0/ra
      -- 
    ra_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_150_load_0_ack_0, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	67 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	28 
    -- CP-element group 19: 	30 
    -- CP-element group 19: 	32 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (33) 
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/$exit
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/merge_req
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/ptr_deref_150_Merge/merge_ack
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/rr
      -- 
    ca_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_150_load_0_ack_1, ack => sendOutput_CP_26_elements(19)); -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_154_inst_req_0); -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_164_inst_req_0); -- 
    rr_391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_174_inst_req_0); -- 
    rr_405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_184_inst_req_0); -- 
    rr_419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_194_inst_req_0); -- 
    rr_433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_204_inst_req_0); -- 
    rr_447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_214_inst_req_0); -- 
    rr_461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(19), ack => type_cast_224_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Sample/ra
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_154_inst_ack_0, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	67 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/ca
      -- 
    ca_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_154_inst_ack_1, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Sample/ra
      -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	67 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	53 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/ca
      -- 
    ca_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Sample/ra
      -- 
    ra_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_174_inst_ack_0, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	67 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/ca
      -- 
    ca_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_174_inst_ack_1, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Sample/ra
      -- 
    ra_406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_184_inst_ack_0, ack => sendOutput_CP_26_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	67 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	47 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/ca
      -- 
    ca_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_184_inst_ack_1, ack => sendOutput_CP_26_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Sample/ra
      -- 
    ra_420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	44 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/ca
      -- 
    ca_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => sendOutput_CP_26_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	19 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Sample/ra
      -- 
    ra_434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_204_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	67 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	41 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/ca
      -- 
    ca_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_204_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	19 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Sample/ra
      -- 
    ra_448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => sendOutput_CP_26_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	67 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/ca
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => sendOutput_CP_26_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	19 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Sample/ra
      -- 
    ra_462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_0, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	67 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/req
      -- 
    ca_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_1, ack => sendOutput_CP_26_elements(35)); -- 
    req_475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_226_inst_req_0); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_update_start_
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/req
      -- 
    ack_476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_226_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_226_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_226_Update/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_226_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/req
      -- 
    req_489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_229_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(33) & sendOutput_CP_26_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_update_start_
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/req
      -- 
    ack_490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_229_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_229_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_229_Update/ack
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_229_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	31 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/req
      -- 
    req_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_232_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(31) & sendOutput_CP_26_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_update_start_
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/req
      -- 
    ack_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_232_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_232_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_232_Update/ack
      -- 
    ack_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_232_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/req
      -- 
    req_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_235_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(29) & sendOutput_CP_26_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_update_start_
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/req
      -- 
    ack_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_235_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_235_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_235_Update/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_235_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	27 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/req
      -- 
    req_531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_238_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(27) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_update_start_
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/req
      -- 
    ack_532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_238_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_238_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_238_Update/ack
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_238_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/req
      -- 
    req_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => WPIPE_zeropad_output_pipe_241_inst_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(25) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_update_start_
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/req
      -- 
    ack_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_241_inst_ack_0, ack => sendOutput_CP_26_elements(51)); -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(51), ack => WPIPE_zeropad_output_pipe_241_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_241_Update/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_241_inst_ack_1, ack => sendOutput_CP_26_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	23 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/req
      -- 
    req_559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => WPIPE_zeropad_output_pipe_244_inst_req_0); -- 
    sendOutput_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(23) & sendOutput_CP_26_elements(52);
      gj_sendOutput_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_update_start_
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/req
      -- 
    ack_560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_244_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(54), ack => WPIPE_zeropad_output_pipe_244_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_244_Update/ack
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_244_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/req
      -- 
    req_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => WPIPE_zeropad_output_pipe_247_inst_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(21) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_update_start_
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/req
      -- 
    ack_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_247_inst_ack_0, ack => sendOutput_CP_26_elements(57)); -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(57), ack => WPIPE_zeropad_output_pipe_247_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/WPIPE_zeropad_output_pipe_247_Update/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_247_inst_ack_1, ack => sendOutput_CP_26_elements(58)); -- 
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260__exit__
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261__entry__
      -- CP-element group 59: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/$exit
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_27/R_exitcond9_262_place
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_27/if_stmt_261_else_link/$entry
      -- 
    branch_req_587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(59), ack => if_stmt_261_branch_req_0); -- 
    sendOutput_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(14) & sendOutput_CP_26_elements(58);
      gj_sendOutput_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  merge  transition  place  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267__exit__
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xendx_xloopexit_forx_xend
      -- CP-element group 60: 	 branch_block_stmt_27/if_stmt_261_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_27/if_stmt_261_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_27/merge_stmt_267_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_27/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_261_branch_ack_1, ack => sendOutput_CP_26_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	64 
    -- CP-element group 61:  members (12) 
      -- CP-element group 61: 	 branch_block_stmt_27/if_stmt_261_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_27/if_stmt_261_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/cr
      -- 
    else_choice_transition_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_261_branch_ack_0, ack => sendOutput_CP_26_elements(61)); -- 
    rr_640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_139_inst_req_0); -- 
    cr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(61), ack => type_cast_139_inst_req_1); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	13 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/$exit
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_137_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_27/bbx_xnph_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_req
      -- 
    phi_stmt_133_req_621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_req_621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(62), ack => phi_stmt_133_req_0); -- 
    -- Element group sendOutput_CP_26_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(13), ack => sendOutput_CP_26_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Sample/ra
      -- 
    ra_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => sendOutput_CP_26_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	61 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/Update/ca
      -- 
    ca_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => sendOutput_CP_26_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_sources/type_cast_139/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_27/forx_xbody_forx_xbody_PhiReq/phi_stmt_133/phi_stmt_133_req
      -- 
    phi_stmt_133_req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(65), ack => phi_stmt_133_req_1); -- 
    sendOutput_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(63) & sendOutput_CP_26_elements(64);
      gj_sendOutput_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_27/merge_stmt_132_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_27/merge_stmt_132_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(66) <= OrReduce(sendOutput_CP_26_elements(62) & sendOutput_CP_26_elements(65));
    -- CP-element group 67:  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: 	15 
    -- CP-element group 67: 	17 
    -- CP-element group 67: 	19 
    -- CP-element group 67: 	21 
    -- CP-element group 67: 	23 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	27 
    -- CP-element group 67: 	29 
    -- CP-element group 67: 	31 
    -- CP-element group 67: 	33 
    -- CP-element group 67: 	35 
    -- CP-element group 67:  members (53) 
      -- CP-element group 67: 	 branch_block_stmt_27/merge_stmt_132__exit__
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260__entry__
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_164_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resized_1
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scaled_1
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_computed_1
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/index_resize_req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_resize_1/index_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/scale_rename_req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_index_scale_1/scale_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_update_start
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/array_obj_ref_145_final_index_sum_regn_Update/req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/addr_of_146_complete/req
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/ptr_deref_150_Update/word_access_complete/word_0/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_154_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_174_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_184_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_194_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_204_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_214_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_update_start_
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_27/assign_stmt_147_to_assign_stmt_260/type_cast_224_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_27/merge_stmt_132_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/merge_stmt_132_PhiAck/phi_stmt_133_ack
      -- 
    phi_stmt_133_ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_133_ack_0, ack => sendOutput_CP_26_elements(67)); -- 
    cr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_164_inst_req_1); -- 
    req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_145_index_offset_req_0); -- 
    req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => array_obj_ref_145_index_offset_req_1); -- 
    req_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => addr_of_146_final_reg_req_1); -- 
    cr_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => ptr_deref_150_load_0_req_1); -- 
    cr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_154_inst_req_1); -- 
    cr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_174_inst_req_1); -- 
    cr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_184_inst_req_1); -- 
    cr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_194_inst_req_1); -- 
    cr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_204_inst_req_1); -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_214_inst_req_1); -- 
    cr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(67), ack => type_cast_224_inst_req_1); -- 
    -- CP-element group 68:  merge  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	10 
    -- CP-element group 68: 	60 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_27/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/branch_block_stmt_27__exit__
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269__exit__
      -- CP-element group 68: 	 branch_block_stmt_27/return__
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271__exit__
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_269_PhiAck/dummy
      -- CP-element group 68: 	 branch_block_stmt_27/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_27/merge_stmt_271_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(68) <= OrReduce(sendOutput_CP_26_elements(10) & sendOutput_CP_26_elements(60));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_144_resized : std_logic_vector(13 downto 0);
    signal R_indvar_144_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_145_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_147 : std_logic_vector(31 downto 0);
    signal cmp77_90 : std_logic_vector(0 downto 0);
    signal conv14_155 : std_logic_vector(7 downto 0);
    signal conv20_165 : std_logic_vector(7 downto 0);
    signal conv26_175 : std_logic_vector(7 downto 0);
    signal conv32_185 : std_logic_vector(7 downto 0);
    signal conv38_195 : std_logic_vector(7 downto 0);
    signal conv44_205 : std_logic_vector(7 downto 0);
    signal conv50_215 : std_logic_vector(7 downto 0);
    signal conv56_225 : std_logic_vector(7 downto 0);
    signal conv_77 : std_logic_vector(63 downto 0);
    signal exitcond9_260 : std_logic_vector(0 downto 0);
    signal iNsTr_0_35 : std_logic_vector(31 downto 0);
    signal iNsTr_1_47 : std_logic_vector(31 downto 0);
    signal iNsTr_2_59 : std_logic_vector(31 downto 0);
    signal indvar_133 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_255 : std_logic_vector(63 downto 0);
    signal mul3_73 : std_logic_vector(31 downto 0);
    signal mul_68 : std_logic_vector(31 downto 0);
    signal ptr_deref_150_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_150_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_150_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_150_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_150_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_38_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_38_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_38_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_38_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_38_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_50_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_50_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_50_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_50_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_50_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_62_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_62_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_62_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_62_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_62_word_offset_0 : std_logic_vector(6 downto 0);
    signal shr17_161 : std_logic_vector(63 downto 0);
    signal shr23_171 : std_logic_vector(63 downto 0);
    signal shr29_181 : std_logic_vector(63 downto 0);
    signal shr35_191 : std_logic_vector(63 downto 0);
    signal shr41_201 : std_logic_vector(63 downto 0);
    signal shr47_211 : std_logic_vector(63 downto 0);
    signal shr53_221 : std_logic_vector(63 downto 0);
    signal shr76x_xmask_83 : std_logic_vector(63 downto 0);
    signal tmp11_151 : std_logic_vector(63 downto 0);
    signal tmp1_51 : std_logic_vector(31 downto 0);
    signal tmp2_63 : std_logic_vector(31 downto 0);
    signal tmp3_102 : std_logic_vector(31 downto 0);
    signal tmp4_107 : std_logic_vector(31 downto 0);
    signal tmp5_111 : std_logic_vector(63 downto 0);
    signal tmp6_117 : std_logic_vector(63 downto 0);
    signal tmp7_123 : std_logic_vector(0 downto 0);
    signal tmp_39 : std_logic_vector(31 downto 0);
    signal type_cast_115_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_121_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_128_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_137_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_139_wire : std_logic_vector(63 downto 0);
    signal type_cast_159_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_179_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_189_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_209_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_253_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_81_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_87_wire_constant : std_logic_vector(63 downto 0);
    signal umax8_130 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_145_constant_part_of_offset <= "00000000000000";
    array_obj_ref_145_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_145_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_145_resized_base_address <= "00000000000000";
    iNsTr_0_35 <= "00000000000000000000000000000011";
    iNsTr_1_47 <= "00000000000000000000000000000100";
    iNsTr_2_59 <= "00000000000000000000000000000101";
    ptr_deref_150_word_offset_0 <= "00000000000000";
    ptr_deref_38_word_offset_0 <= "0000000";
    ptr_deref_50_word_offset_0 <= "0000000";
    ptr_deref_62_word_offset_0 <= "0000000";
    type_cast_115_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_121_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_128_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_137_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_159_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_179_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_189_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_199_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_209_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_253_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_81_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_87_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_133: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_137_wire_constant & type_cast_139_wire;
      req <= phi_stmt_133_req_0 & phi_stmt_133_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_133",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_133_ack_0,
          idata => idata,
          odata => indvar_133,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_133
    -- flow-through select operator MUX_129_inst
    umax8_130 <= tmp6_117 when (tmp7_123(0) /=  '0') else type_cast_128_wire_constant;
    addr_of_146_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_146_final_reg_req_0;
      addr_of_146_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_146_final_reg_req_1;
      addr_of_146_final_reg_ack_1<= rack(0);
      addr_of_146_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_146_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_145_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_110_inst_req_0;
      type_cast_110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_110_inst_req_1;
      type_cast_110_inst_ack_1<= rack(0);
      type_cast_110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_139_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_154_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_154_inst_req_0;
      type_cast_154_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_154_inst_req_1;
      type_cast_154_inst_ack_1<= rack(0);
      type_cast_154_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_154_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_155,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_174_inst_req_0;
      type_cast_174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_174_inst_req_1;
      type_cast_174_inst_ack_1<= rack(0);
      type_cast_174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_184_inst_req_0;
      type_cast_184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_184_inst_req_1;
      type_cast_184_inst_ack_1<= rack(0);
      type_cast_184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_181,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_185,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_204_inst_req_0;
      type_cast_204_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_204_inst_req_1;
      type_cast_204_inst_ack_1<= rack(0);
      type_cast_204_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_205,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_224_inst_req_0;
      type_cast_224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_224_inst_req_1;
      type_cast_224_inst_ack_1<= rack(0);
      type_cast_224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr53_221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul3_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_145_index_1_rename
    process(R_indvar_144_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_144_resized;
      ov(13 downto 0) := iv;
      R_indvar_144_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_145_index_1_resize
    process(indvar_133) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_133;
      ov := iv(13 downto 0);
      R_indvar_144_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_145_root_address_inst
    process(array_obj_ref_145_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_145_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_145_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_addr_0
    process(ptr_deref_150_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_150_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_150_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_base_resize
    process(arrayidx_147) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_147;
      ov := iv(13 downto 0);
      ptr_deref_150_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_gather_scatter
    process(ptr_deref_150_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_150_data_0;
      ov(63 downto 0) := iv;
      tmp11_151 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_150_root_address_inst
    process(ptr_deref_150_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_150_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_150_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_addr_0
    process(ptr_deref_38_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_38_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_38_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_base_resize
    process(iNsTr_0_35) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_35;
      ov := iv(6 downto 0);
      ptr_deref_38_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_gather_scatter
    process(ptr_deref_38_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_38_data_0;
      ov(31 downto 0) := iv;
      tmp_39 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_38_root_address_inst
    process(ptr_deref_38_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_38_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_38_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_addr_0
    process(ptr_deref_50_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_50_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_50_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_base_resize
    process(iNsTr_1_47) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_47;
      ov := iv(6 downto 0);
      ptr_deref_50_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_gather_scatter
    process(ptr_deref_50_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_50_data_0;
      ov(31 downto 0) := iv;
      tmp1_51 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_50_root_address_inst
    process(ptr_deref_50_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_50_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_50_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_addr_0
    process(ptr_deref_62_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_62_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_62_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_base_resize
    process(iNsTr_2_59) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_59;
      ov := iv(6 downto 0);
      ptr_deref_62_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_gather_scatter
    process(ptr_deref_62_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_62_data_0;
      ov(31 downto 0) := iv;
      tmp2_63 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_62_root_address_inst
    process(ptr_deref_62_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_62_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_62_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_261_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_260;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_261_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_261_branch_req_0,
          ack0 => if_stmt_261_branch_ack_0,
          ack1 => if_stmt_261_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_91_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_90;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_91_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_91_branch_req_0,
          ack0 => if_stmt_91_branch_ack_0,
          ack1 => if_stmt_91_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_254_inst
    process(indvar_133) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_133, type_cast_253_wire_constant, tmp_var);
      indvarx_xnext_255 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_82_inst
    process(conv_77) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv_77, type_cast_81_wire_constant, tmp_var);
      shr76x_xmask_83 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_259_inst
    process(indvarx_xnext_255, umax8_130) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_255, umax8_130, tmp_var);
      exitcond9_260 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_88_inst
    process(shr76x_xmask_83) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr76x_xmask_83, type_cast_87_wire_constant, tmp_var);
      cmp77_90 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_116_inst
    process(tmp5_111) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_111, type_cast_115_wire_constant, tmp_var);
      tmp6_117 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_160_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_159_wire_constant, tmp_var);
      shr17_161 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_170_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_169_wire_constant, tmp_var);
      shr23_171 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_180_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_179_wire_constant, tmp_var);
      shr29_181 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_190_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_189_wire_constant, tmp_var);
      shr35_191 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_200_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_199_wire_constant, tmp_var);
      shr41_201 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_210_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_209_wire_constant, tmp_var);
      shr47_211 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_220_inst
    process(tmp11_151) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp11_151, type_cast_219_wire_constant, tmp_var);
      shr53_221 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_101_inst
    process(tmp1_51, tmp_39) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_51, tmp_39, tmp_var);
      tmp3_102 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_106_inst
    process(tmp3_102, tmp2_63) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_102, tmp2_63, tmp_var);
      tmp4_107 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_67_inst
    process(tmp1_51, tmp_39) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_51, tmp_39, tmp_var);
      mul_68 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_72_inst
    process(mul_68, tmp2_63) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_68, tmp2_63, tmp_var);
      mul3_73 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_122_inst
    process(tmp6_117) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp6_117, type_cast_121_wire_constant, tmp_var);
      tmp7_123 <= tmp_var; --
    end process;
    -- shared split operator group (17) : array_obj_ref_145_index_offset 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_144_scaled;
      array_obj_ref_145_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_145_index_offset_req_0;
      array_obj_ref_145_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_145_index_offset_req_1;
      array_obj_ref_145_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_17_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared load operator group (0) : ptr_deref_150_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_150_load_0_req_0;
      ptr_deref_150_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_150_load_0_req_1;
      ptr_deref_150_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_150_word_address_0;
      ptr_deref_150_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_38_load_0 ptr_deref_50_load_0 ptr_deref_62_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_38_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_50_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_62_load_0_req_0;
      ptr_deref_38_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_50_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_62_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_38_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_50_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_62_load_0_req_1;
      ptr_deref_38_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_50_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_62_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_38_word_address_0 & ptr_deref_50_word_address_0 & ptr_deref_62_word_address_0;
      ptr_deref_38_data_0 <= data_out(95 downto 64);
      ptr_deref_50_data_0 <= data_out(63 downto 32);
      ptr_deref_62_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(6 downto 0),
          mtag => memory_space_6_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_226_inst WPIPE_zeropad_output_pipe_229_inst WPIPE_zeropad_output_pipe_232_inst WPIPE_zeropad_output_pipe_235_inst WPIPE_zeropad_output_pipe_238_inst WPIPE_zeropad_output_pipe_241_inst WPIPE_zeropad_output_pipe_244_inst WPIPE_zeropad_output_pipe_247_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_226_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_229_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_232_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_235_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_238_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_241_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_244_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_247_inst_req_0;
      WPIPE_zeropad_output_pipe_226_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_229_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_232_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_235_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_238_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_241_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_244_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_247_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_226_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_229_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_232_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_235_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_238_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_241_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_244_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_247_inst_req_1;
      WPIPE_zeropad_output_pipe_226_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_229_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_232_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_235_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_238_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_241_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_244_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_247_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv56_225 & conv50_215 & conv44_205 & conv38_195 & conv32_185 & conv26_175 & conv20_165 & conv14_155;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_684_start: Boolean;
  signal testConfigure_CP_684_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal STORE_row_high_326_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_ack_1 : boolean;
  signal type_cast_595_inst_req_1 : boolean;
  signal type_cast_595_inst_ack_0 : boolean;
  signal type_cast_595_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_req_1 : boolean;
  signal ptr_deref_320_store_0_ack_0 : boolean;
  signal type_cast_595_inst_ack_1 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_330_inst_ack_0 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_req_0 : boolean;
  signal STORE_row_high_326_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_ack_0 : boolean;
  signal STORE_row_high_326_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_307_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_ack_0 : boolean;
  signal type_cast_294_inst_ack_1 : boolean;
  signal type_cast_294_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_req_0 : boolean;
  signal type_cast_294_inst_ack_0 : boolean;
  signal type_cast_294_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_ack_1 : boolean;
  signal type_cast_311_inst_ack_1 : boolean;
  signal type_cast_311_inst_req_1 : boolean;
  signal ptr_deref_285_store_0_ack_1 : boolean;
  signal ptr_deref_303_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_req_0 : boolean;
  signal ptr_deref_285_store_0_req_1 : boolean;
  signal ptr_deref_303_store_0_req_1 : boolean;
  signal type_cast_613_inst_req_0 : boolean;
  signal type_cast_528_inst_req_1 : boolean;
  signal ptr_deref_320_store_0_req_0 : boolean;
  signal ptr_deref_303_store_0_ack_0 : boolean;
  signal ptr_deref_285_store_0_ack_0 : boolean;
  signal type_cast_613_inst_ack_0 : boolean;
  signal ptr_deref_285_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_609_inst_ack_0 : boolean;
  signal ptr_deref_303_store_0_req_0 : boolean;
  signal type_cast_631_inst_req_0 : boolean;
  signal type_cast_682_inst_req_0 : boolean;
  signal type_cast_682_inst_ack_1 : boolean;
  signal phi_stmt_508_req_0 : boolean;
  signal array_obj_ref_520_index_offset_req_0 : boolean;
  signal type_cast_311_inst_ack_0 : boolean;
  signal type_cast_311_inst_req_0 : boolean;
  signal ptr_deref_320_store_0_ack_1 : boolean;
  signal ptr_deref_320_store_0_req_1 : boolean;
  signal type_cast_631_inst_ack_0 : boolean;
  signal type_cast_528_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_ack_1 : boolean;
  signal STORE_row_high_326_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_324_inst_req_1 : boolean;
  signal array_obj_ref_520_index_offset_ack_0 : boolean;
  signal type_cast_613_inst_req_1 : boolean;
  signal type_cast_613_inst_ack_1 : boolean;
  signal addr_of_521_final_reg_req_0 : boolean;
  signal addr_of_521_final_reg_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_req_0 : boolean;
  signal type_cast_631_inst_req_1 : boolean;
  signal type_cast_631_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_req_0 : boolean;
  signal addr_of_521_final_reg_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_ack_0 : boolean;
  signal addr_of_521_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_req_1 : boolean;
  signal type_cast_514_inst_ack_1 : boolean;
  signal if_stmt_671_branch_req_0 : boolean;
  signal phi_stmt_508_req_1 : boolean;
  signal type_cast_514_inst_req_1 : boolean;
  signal type_cast_514_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_537_inst_ack_1 : boolean;
  signal type_cast_514_inst_ack_0 : boolean;
  signal array_obj_ref_520_index_offset_req_1 : boolean;
  signal array_obj_ref_520_index_offset_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_627_inst_ack_1 : boolean;
  signal type_cast_682_inst_req_1 : boolean;
  signal type_cast_541_inst_req_0 : boolean;
  signal type_cast_541_inst_ack_0 : boolean;
  signal type_cast_541_inst_req_1 : boolean;
  signal if_stmt_671_branch_ack_0 : boolean;
  signal type_cast_682_inst_ack_0 : boolean;
  signal type_cast_541_inst_ack_1 : boolean;
  signal type_cast_559_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_290_inst_ack_1 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_req_1 : boolean;
  signal STORE_col_high_332_store_0_req_0 : boolean;
  signal STORE_col_high_332_store_0_ack_0 : boolean;
  signal STORE_col_high_332_store_0_req_1 : boolean;
  signal STORE_col_high_332_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_336_inst_ack_1 : boolean;
  signal ptr_deref_657_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_req_1 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal STORE_depth_high_338_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_ack_0 : boolean;
  signal STORE_depth_high_338_store_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_ack_0 : boolean;
  signal STORE_depth_high_338_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_591_inst_req_0 : boolean;
  signal STORE_depth_high_338_store_0_ack_1 : boolean;
  signal ptr_deref_657_store_0_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_req_1 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_342_inst_ack_1 : boolean;
  signal if_stmt_671_branch_ack_1 : boolean;
  signal type_cast_577_inst_ack_1 : boolean;
  signal type_cast_577_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_555_inst_req_0 : boolean;
  signal STORE_pad_344_store_0_req_0 : boolean;
  signal STORE_pad_344_store_0_ack_0 : boolean;
  signal STORE_pad_344_store_0_req_1 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal STORE_pad_344_store_0_ack_1 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_348_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_req_1 : boolean;
  signal type_cast_352_inst_req_0 : boolean;
  signal type_cast_352_inst_ack_0 : boolean;
  signal type_cast_352_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_ack_1 : boolean;
  signal type_cast_352_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_573_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_524_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_ack_0 : boolean;
  signal ptr_deref_363_store_0_req_0 : boolean;
  signal ptr_deref_363_store_0_ack_0 : boolean;
  signal ptr_deref_363_store_0_req_1 : boolean;
  signal ptr_deref_363_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_645_inst_req_0 : boolean;
  signal type_cast_559_inst_ack_1 : boolean;
  signal type_cast_559_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_1 : boolean;
  signal ptr_deref_657_store_0_ack_0 : boolean;
  signal type_cast_559_inst_ack_0 : boolean;
  signal ptr_deref_657_store_0_req_0 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal ptr_deref_382_store_0_req_0 : boolean;
  signal ptr_deref_382_store_0_ack_0 : boolean;
  signal ptr_deref_382_store_0_req_1 : boolean;
  signal ptr_deref_382_store_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_386_inst_ack_1 : boolean;
  signal type_cast_390_inst_req_0 : boolean;
  signal type_cast_390_inst_ack_0 : boolean;
  signal type_cast_390_inst_req_1 : boolean;
  signal type_cast_390_inst_ack_1 : boolean;
  signal ptr_deref_401_store_0_req_0 : boolean;
  signal ptr_deref_401_store_0_ack_0 : boolean;
  signal ptr_deref_401_store_0_req_1 : boolean;
  signal ptr_deref_401_store_0_ack_1 : boolean;
  signal ptr_deref_414_load_0_req_0 : boolean;
  signal ptr_deref_414_load_0_ack_0 : boolean;
  signal ptr_deref_414_load_0_req_1 : boolean;
  signal ptr_deref_414_load_0_ack_1 : boolean;
  signal ptr_deref_426_load_0_req_0 : boolean;
  signal ptr_deref_426_load_0_ack_0 : boolean;
  signal ptr_deref_426_load_0_req_1 : boolean;
  signal ptr_deref_426_load_0_ack_1 : boolean;
  signal ptr_deref_438_load_0_req_0 : boolean;
  signal ptr_deref_438_load_0_ack_0 : boolean;
  signal ptr_deref_438_load_0_req_1 : boolean;
  signal ptr_deref_438_load_0_ack_1 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal if_stmt_466_branch_req_0 : boolean;
  signal if_stmt_466_branch_ack_1 : boolean;
  signal if_stmt_466_branch_ack_0 : boolean;
  signal type_cast_485_inst_req_0 : boolean;
  signal type_cast_485_inst_ack_0 : boolean;
  signal type_cast_485_inst_req_1 : boolean;
  signal type_cast_485_inst_ack_1 : boolean;
  signal phi_stmt_508_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_684_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_684_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_684: Block -- control-path 
    signal testConfigure_CP_684_elements: BooleanArray(132 downto 0);
    -- 
  begin -- 
    testConfigure_CP_684_elements(0) <= testConfigure_CP_684_start;
    testConfigure_CP_684_symbol <= testConfigure_CP_684_elements(125);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	14 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	50 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0:  members (252) 
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465__entry__
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/branch_block_stmt_277__entry__
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/split_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/split_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/ptr_deref_285_Split/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_address_resized
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_update_start_
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/cr
      -- 
    cr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_row_high_326_store_0_req_1); -- 
    cr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_294_inst_req_1); -- 
    rr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => RPIPE_zeropad_input_pipe_290_inst_req_0); -- 
    cr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_311_inst_req_1); -- 
    cr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_285_store_0_req_1); -- 
    cr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_303_store_0_req_1); -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_285_store_0_req_0); -- 
    cr_921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_320_store_0_req_1); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_col_high_332_store_0_req_1); -- 
    cr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_depth_high_338_store_0_req_1); -- 
    cr_1109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => STORE_pad_344_store_0_req_1); -- 
    cr_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_352_inst_req_1); -- 
    cr_1187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_363_store_0_req_1); -- 
    cr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_371_inst_req_1); -- 
    cr_1265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_382_store_0_req_1); -- 
    cr_1293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_390_inst_req_1); -- 
    cr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_401_store_0_req_1); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_414_load_0_req_1); -- 
    cr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_426_load_0_req_1); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => ptr_deref_438_load_0_req_1); -- 
    cr_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(0), ack => type_cast_452_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	70 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Sample/$exit
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_285_store_0_ack_0, ack => testConfigure_CP_684_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	77 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_update_completed_
      -- 
    ca_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_285_store_0_ack_1, ack => testConfigure_CP_684_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_update_start_
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_sample_completed_
      -- 
    ra_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_290_inst_ack_0, ack => testConfigure_CP_684_elements(3)); -- 
    cr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(3), ack => RPIPE_zeropad_input_pipe_290_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_290_Update/ca
      -- 
    ca_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_290_inst_ack_1, ack => testConfigure_CP_684_elements(4)); -- 
    rr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(4), ack => type_cast_294_inst_req_0); -- 
    rr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(4), ack => RPIPE_zeropad_input_pipe_307_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_sample_completed_
      -- 
    ra_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_294_inst_ack_0, ack => testConfigure_CP_684_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_294_update_completed_
      -- 
    ca_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_294_inst_ack_1, ack => testConfigure_CP_684_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	70 
    -- CP-element group 7: 	0 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/rr
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/split_ack
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/split_req
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/$exit
      -- CP-element group 7: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/ptr_deref_303_Split/$entry
      -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(7), ack => ptr_deref_303_store_0_req_0); -- 
    testConfigure_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(70) & testConfigure_CP_684_elements(0) & testConfigure_CP_684_elements(6);
      gj_testConfigure_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/ra
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Sample/word_access_start/$exit
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_303_store_0_ack_0, ack => testConfigure_CP_684_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	77 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_update_completed_
      -- 
    ca_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_303_store_0_ack_1, ack => testConfigure_CP_684_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_update_start_
      -- CP-element group 10: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_sample_completed_
      -- 
    ra_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_307_inst_ack_0, ack => testConfigure_CP_684_elements(10)); -- 
    cr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(10), ack => RPIPE_zeropad_input_pipe_307_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_307_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_sample_start_
      -- 
    ca_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_307_inst_ack_1, ack => testConfigure_CP_684_elements(11)); -- 
    rr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(11), ack => type_cast_311_inst_req_0); -- 
    rr_930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(11), ack => RPIPE_zeropad_input_pipe_324_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_sample_completed_
      -- 
    ra_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_0, ack => testConfigure_CP_684_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_311_update_completed_
      -- 
    ca_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_1, ack => testConfigure_CP_684_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: 	71 
    -- CP-element group 14: 	0 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/rr
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/split_ack
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/split_req
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/$exit
      -- CP-element group 14: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/ptr_deref_320_Split/$entry
      -- 
    rr_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(14), ack => ptr_deref_320_store_0_req_0); -- 
    testConfigure_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(13) & testConfigure_CP_684_elements(71) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	72 
    -- CP-element group 15: 	73 
    -- CP-element group 15: 	74 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Sample/$exit
      -- 
    ra_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_store_0_ack_0, ack => testConfigure_CP_684_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	77 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_Update/word_access_complete/word_0/ca
      -- 
    ca_922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_store_0_ack_1, ack => testConfigure_CP_684_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_update_start_
      -- CP-element group 17: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/cr
      -- 
    ra_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_324_inst_ack_0, ack => testConfigure_CP_684_elements(17)); -- 
    cr_935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(17), ack => RPIPE_zeropad_input_pipe_324_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_324_Update/ca
      -- 
    ca_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_324_inst_ack_1, ack => testConfigure_CP_684_elements(18)); -- 
    rr_977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(18), ack => RPIPE_zeropad_input_pipe_330_inst_req_0); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/rr
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/split_ack
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/split_req
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/$exit
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/STORE_row_high_326_Split/$entry
      -- CP-element group 19: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/$entry
      -- 
    rr_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(19), ack => STORE_row_high_326_store_0_req_0); -- 
    testConfigure_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(18) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/ra
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Sample/$exit
      -- 
    ra_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_326_store_0_ack_0, ack => testConfigure_CP_684_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	77 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_row_high_326_Update/word_access_complete/word_0/ca
      -- 
    ca_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_326_store_0_ack_1, ack => testConfigure_CP_684_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_update_start_
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Sample/ra
      -- 
    ra_978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_330_inst_ack_0, ack => testConfigure_CP_684_elements(22)); -- 
    cr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(22), ack => RPIPE_zeropad_input_pipe_330_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	27 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_330_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/rr
      -- 
    ca_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_330_inst_ack_1, ack => testConfigure_CP_684_elements(23)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(23), ack => RPIPE_zeropad_input_pipe_336_inst_req_0); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/$exit
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/split_req
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/STORE_col_high_332_Split/split_ack
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/rr
      -- 
    rr_1004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(24), ack => STORE_col_high_332_store_0_req_0); -- 
    testConfigure_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(23) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Sample/word_access_start/word_0/ra
      -- 
    ra_1005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_332_store_0_ack_0, ack => testConfigure_CP_684_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	77 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_col_high_332_Update/word_access_complete/word_0/ca
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_332_store_0_ack_1, ack => testConfigure_CP_684_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_update_start_
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/cr
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_336_inst_ack_0, ack => testConfigure_CP_684_elements(27)); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(27), ack => RPIPE_zeropad_input_pipe_336_inst_req_1); -- 
    -- CP-element group 28:  fork  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	32 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_336_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/rr
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_336_inst_ack_1, ack => testConfigure_CP_684_elements(28)); -- 
    rr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(28), ack => RPIPE_zeropad_input_pipe_342_inst_req_0); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/$exit
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/split_req
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/STORE_depth_high_338_Split/split_ack
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/rr
      -- 
    rr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(29), ack => STORE_depth_high_338_store_0_req_0); -- 
    testConfigure_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(28) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Sample/word_access_start/word_0/ra
      -- 
    ra_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_338_store_0_ack_0, ack => testConfigure_CP_684_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	77 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_depth_high_338_Update/word_access_complete/word_0/ca
      -- 
    ca_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_338_store_0_ack_1, ack => testConfigure_CP_684_elements(31)); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	28 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_update_start_
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/cr
      -- 
    ra_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_342_inst_ack_0, ack => testConfigure_CP_684_elements(32)); -- 
    cr_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(32), ack => RPIPE_zeropad_input_pipe_342_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	37 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_342_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/rr
      -- 
    ca_1077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_342_inst_ack_1, ack => testConfigure_CP_684_elements(33)); -- 
    rr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(33), ack => RPIPE_zeropad_input_pipe_348_inst_req_0); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/$exit
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/split_req
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/STORE_pad_344_Split/split_ack
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/rr
      -- 
    rr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(34), ack => STORE_pad_344_store_0_req_0); -- 
    testConfigure_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(33) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Sample/word_access_start/word_0/ra
      -- 
    ra_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_344_store_0_ack_0, ack => testConfigure_CP_684_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	77 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/STORE_pad_344_Update/word_access_complete/word_0/ca
      -- 
    ca_1110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_344_store_0_ack_1, ack => testConfigure_CP_684_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	33 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_update_start_
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/cr
      -- 
    ra_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_348_inst_ack_0, ack => testConfigure_CP_684_elements(37)); -- 
    cr_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(37), ack => RPIPE_zeropad_input_pipe_348_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	44 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_348_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/rr
      -- 
    ca_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_348_inst_ack_1, ack => testConfigure_CP_684_elements(38)); -- 
    rr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(38), ack => type_cast_352_inst_req_0); -- 
    rr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(38), ack => RPIPE_zeropad_input_pipe_367_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Sample/ra
      -- 
    ra_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_0, ack => testConfigure_CP_684_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_352_Update/ca
      -- 
    ca_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_1, ack => testConfigure_CP_684_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/$exit
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/split_req
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/ptr_deref_363_Split/split_ack
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/rr
      -- 
    rr_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(41), ack => ptr_deref_363_store_0_req_0); -- 
    testConfigure_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(40) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	75 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Sample/word_access_start/word_0/ra
      -- 
    ra_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_store_0_ack_0, ack => testConfigure_CP_684_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	77 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_Update/word_access_complete/word_0/ca
      -- 
    ca_1188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_store_0_ack_1, ack => testConfigure_CP_684_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	38 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_update_start_
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/cr
      -- 
    ra_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_0, ack => testConfigure_CP_684_elements(44)); -- 
    cr_1201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(44), ack => RPIPE_zeropad_input_pipe_367_inst_req_1); -- 
    -- CP-element group 45:  fork  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	51 
    -- CP-element group 45:  members (9) 
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_367_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/rr
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/rr
      -- 
    ca_1202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_1, ack => testConfigure_CP_684_elements(45)); -- 
    rr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(45), ack => type_cast_371_inst_req_0); -- 
    rr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(45), ack => RPIPE_zeropad_input_pipe_386_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Sample/ra
      -- 
    ra_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => testConfigure_CP_684_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_371_Update/ca
      -- 
    ca_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => testConfigure_CP_684_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	75 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/ptr_deref_382_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/rr
      -- 
    rr_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(48), ack => ptr_deref_382_store_0_req_0); -- 
    testConfigure_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(47) & testConfigure_CP_684_elements(75) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	76 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Sample/word_access_start/word_0/ra
      -- 
    ra_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_382_store_0_ack_0, ack => testConfigure_CP_684_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	0 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	77 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_Update/word_access_complete/word_0/ca
      -- 
    ca_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_382_store_0_ack_1, ack => testConfigure_CP_684_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	45 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_update_start_
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/cr
      -- 
    ra_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_386_inst_ack_0, ack => testConfigure_CP_684_elements(51)); -- 
    cr_1279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(51), ack => RPIPE_zeropad_input_pipe_386_inst_req_1); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/RPIPE_zeropad_input_pipe_386_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/rr
      -- 
    ca_1280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_386_inst_ack_1, ack => testConfigure_CP_684_elements(52)); -- 
    rr_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(52), ack => type_cast_390_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Sample/ra
      -- 
    ra_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_0, ack => testConfigure_CP_684_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_390_Update/ca
      -- 
    ca_1294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_390_inst_ack_1, ack => testConfigure_CP_684_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	76 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/ptr_deref_401_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/rr
      -- 
    rr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(55), ack => ptr_deref_401_store_0_req_0); -- 
    testConfigure_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(54) & testConfigure_CP_684_elements(76) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Sample/word_access_start/word_0/ra
      -- 
    ra_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_401_store_0_ack_0, ack => testConfigure_CP_684_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	77 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_401_Update/word_access_complete/word_0/ca
      -- 
    ca_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_401_store_0_ack_1, ack => testConfigure_CP_684_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	72 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/rr
      -- 
    rr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(58), ack => ptr_deref_414_load_0_req_0); -- 
    testConfigure_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(72) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Sample/word_access_start/word_0/ra
      -- 
    ra_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_414_load_0_ack_0, ack => testConfigure_CP_684_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	67 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_414_Update/ptr_deref_414_Merge/merge_ack
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_414_load_0_ack_1, ack => testConfigure_CP_684_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	73 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/rr
      -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(61), ack => ptr_deref_426_load_0_req_0); -- 
    testConfigure_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(73) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Sample/word_access_start/word_0/ra
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_0, ack => testConfigure_CP_684_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	67 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/word_access_complete/word_0/ca
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/$entry
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/merge_req
      -- CP-element group 63: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_426_Update/ptr_deref_426_Merge/merge_ack
      -- 
    ca_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_1, ack => testConfigure_CP_684_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	74 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/$entry
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/$entry
      -- CP-element group 64: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/rr
      -- 
    rr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(64), ack => ptr_deref_438_load_0_req_0); -- 
    testConfigure_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(74) & testConfigure_CP_684_elements(0);
      gj_testConfigure_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Sample/word_access_start/word_0/ra
      -- 
    ra_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_438_load_0_ack_0, ack => testConfigure_CP_684_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/word_access_complete/word_0/ca
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/$entry
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/$exit
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/merge_req
      -- CP-element group 66: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_438_Update/ptr_deref_438_Merge/merge_ack
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_438_load_0_ack_1, ack => testConfigure_CP_684_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	60 
    -- CP-element group 67: 	63 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/rr
      -- 
    rr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(67), ack => type_cast_452_inst_req_0); -- 
    testConfigure_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(60) & testConfigure_CP_684_elements(63) & testConfigure_CP_684_elements(66);
      gj_testConfigure_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Sample/ra
      -- 
    ra_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => testConfigure_CP_684_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	77 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/type_cast_452_Update/ca
      -- 
    ca_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => testConfigure_CP_684_elements(69)); -- 
    -- CP-element group 70:  transition  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	1 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	7 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_285_ptr_deref_303_delay
      -- 
    -- Element group testConfigure_CP_684_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(1), ack => testConfigure_CP_684_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	8 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	14 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_303_ptr_deref_320_delay
      -- 
    -- Element group testConfigure_CP_684_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(8), ack => testConfigure_CP_684_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  delay-element  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	15 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	58 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_ptr_deref_414_delay
      -- 
    -- Element group testConfigure_CP_684_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(15), ack => testConfigure_CP_684_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  transition  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	15 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	61 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_ptr_deref_426_delay
      -- 
    -- Element group testConfigure_CP_684_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(15), ack => testConfigure_CP_684_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  delay-element  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	15 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	64 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_320_ptr_deref_438_delay
      -- 
    -- Element group testConfigure_CP_684_elements(74) is a control-delay.
    cp_element_74_delay: control_delay_element  generic map(name => " 74_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(15), ack => testConfigure_CP_684_elements(74), clk => clk, reset =>reset);
    -- CP-element group 75:  transition  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	42 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	48 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_363_ptr_deref_382_delay
      -- 
    -- Element group testConfigure_CP_684_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(42), ack => testConfigure_CP_684_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	49 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	55 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/ptr_deref_382_ptr_deref_401_delay
      -- 
    -- Element group testConfigure_CP_684_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(49), ack => testConfigure_CP_684_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  branch  join  transition  place  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	16 
    -- CP-element group 77: 	21 
    -- CP-element group 77: 	26 
    -- CP-element group 77: 	31 
    -- CP-element group 77: 	36 
    -- CP-element group 77: 	43 
    -- CP-element group 77: 	50 
    -- CP-element group 77: 	57 
    -- CP-element group 77: 	69 
    -- CP-element group 77: 	2 
    -- CP-element group 77: 	9 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (10) 
      -- CP-element group 77: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465__exit__
      -- CP-element group 77: 	 branch_block_stmt_277/assign_stmt_283_to_assign_stmt_465/$exit
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466__entry__
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_dead_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_eval_test/$entry
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_eval_test/$exit
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_eval_test/branch_req
      -- CP-element group 77: 	 branch_block_stmt_277/R_cmp71_467_place
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_if_link/$entry
      -- CP-element group 77: 	 branch_block_stmt_277/if_stmt_466_else_link/$entry
      -- 
    branch_req_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(77), ack => if_stmt_466_branch_req_0); -- 
    testConfigure_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(16) & testConfigure_CP_684_elements(21) & testConfigure_CP_684_elements(26) & testConfigure_CP_684_elements(31) & testConfigure_CP_684_elements(36) & testConfigure_CP_684_elements(43) & testConfigure_CP_684_elements(50) & testConfigure_CP_684_elements(57) & testConfigure_CP_684_elements(69) & testConfigure_CP_684_elements(2) & testConfigure_CP_684_elements(9);
      gj_testConfigure_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	132 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_277/if_stmt_466_if_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_277/if_stmt_466_if_link/if_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_277/entry_forx_xend
      -- CP-element group 78: 	 branch_block_stmt_277/entry_forx_xend_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_277/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_466_branch_ack_1, ack => testConfigure_CP_684_elements(78)); -- 
    -- CP-element group 79:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (18) 
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505__entry__
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472__exit__
      -- CP-element group 79: 	 branch_block_stmt_277/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiAck/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_277/merge_stmt_472_PhiAck/dummy
      -- CP-element group 79: 	 branch_block_stmt_277/if_stmt_466_else_link/$exit
      -- CP-element group 79: 	 branch_block_stmt_277/if_stmt_466_else_link/else_choice_transition
      -- CP-element group 79: 	 branch_block_stmt_277/entry_bbx_xnph
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_update_start_
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/cr
      -- 
    else_choice_transition_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_466_branch_ack_0, ack => testConfigure_CP_684_elements(79)); -- 
    rr_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(79), ack => type_cast_485_inst_req_0); -- 
    cr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(79), ack => type_cast_485_inst_req_1); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Sample/ra
      -- 
    ra_1546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_0, ack => testConfigure_CP_684_elements(80)); -- 
    -- CP-element group 81:  transition  place  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	126 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505__exit__
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$entry
      -- CP-element group 81: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/$entry
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/$exit
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_277/assign_stmt_477_to_assign_stmt_505/type_cast_485_Update/ca
      -- 
    ca_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_1, ack => testConfigure_CP_684_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	131 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	121 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_sample_complete
      -- CP-element group 82: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/ack
      -- 
    ack_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_520_index_offset_ack_0, ack => testConfigure_CP_684_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	131 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (11) 
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/$entry
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/$entry
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/req
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/ack
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/$exit
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/sum_rename_req
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_base_plus_offset/sum_rename_ack
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_root_address_calculated
      -- CP-element group 83: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_offset_calculated
      -- 
    ack_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_520_index_offset_ack_1, ack => testConfigure_CP_684_elements(83)); -- 
    req_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(83), ack => addr_of_521_final_reg_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/$exit
      -- CP-element group 84: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_request/ack
      -- CP-element group 84: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_sample_completed_
      -- 
    ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_521_final_reg_ack_0, ack => testConfigure_CP_684_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	131 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (19) 
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/$entry
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/$entry
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_address_resized
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/sum_rename_ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/root_register_req
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_addrgen/root_register_ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/base_resize_req
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_addr_resize/base_resize_ack
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/sum_rename_req
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/$exit
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_plus_offset/$entry
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_root_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_word_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_base_address_calculated
      -- CP-element group 85: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_update_completed_
      -- 
    ack_1600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_521_final_reg_ack_1, ack => testConfigure_CP_684_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	131 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_update_start_
      -- 
    ra_1609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_524_inst_ack_0, ack => testConfigure_CP_684_elements(86)); -- 
    cr_1613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(86), ack => RPIPE_zeropad_input_pipe_524_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_update_completed_
      -- 
    ca_1614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_524_inst_ack_1, ack => testConfigure_CP_684_elements(87)); -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(87), ack => type_cast_528_inst_req_0); -- 
    rr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(87), ack => RPIPE_zeropad_input_pipe_537_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_sample_completed_
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_0, ack => testConfigure_CP_684_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	131 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_update_completed_
      -- 
    ca_1628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_1, ack => testConfigure_CP_684_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_update_start_
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/cr
      -- 
    ra_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_537_inst_ack_0, ack => testConfigure_CP_684_elements(90)); -- 
    cr_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(90), ack => RPIPE_zeropad_input_pipe_537_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_537_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/$entry
      -- 
    ca_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_537_inst_ack_1, ack => testConfigure_CP_684_elements(91)); -- 
    rr_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(91), ack => type_cast_541_inst_req_0); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(91), ack => RPIPE_zeropad_input_pipe_555_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Sample/ra
      -- 
    ra_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_0, ack => testConfigure_CP_684_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	131 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/ca
      -- 
    ca_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_1, ack => testConfigure_CP_684_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_update_start_
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_555_inst_ack_0, ack => testConfigure_CP_684_elements(94)); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(94), ack => RPIPE_zeropad_input_pipe_555_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_555_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_sample_start_
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_555_inst_ack_1, ack => testConfigure_CP_684_elements(95)); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(95), ack => type_cast_559_inst_req_0); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(95), ack => RPIPE_zeropad_input_pipe_573_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_0, ack => testConfigure_CP_684_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	131 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/$exit
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_1, ack => testConfigure_CP_684_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_update_start_
      -- CP-element group 98: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_sample_completed_
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_573_inst_ack_0, ack => testConfigure_CP_684_elements(98)); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(98), ack => RPIPE_zeropad_input_pipe_573_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_573_update_completed_
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_573_inst_ack_1, ack => testConfigure_CP_684_elements(99)); -- 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(99), ack => type_cast_577_inst_req_0); -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(99), ack => RPIPE_zeropad_input_pipe_591_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_sample_completed_
      -- 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => testConfigure_CP_684_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	131 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_update_completed_
      -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_1, ack => testConfigure_CP_684_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_update_start_
      -- CP-element group 102: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_sample_completed_
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_591_inst_ack_0, ack => testConfigure_CP_684_elements(102)); -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(102), ack => RPIPE_zeropad_input_pipe_591_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_591_update_completed_
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_591_inst_ack_1, ack => testConfigure_CP_684_elements(103)); -- 
    rr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(103), ack => type_cast_595_inst_req_0); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(103), ack => RPIPE_zeropad_input_pipe_609_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_sample_completed_
      -- 
    ra_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_0, ack => testConfigure_CP_684_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	131 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_update_completed_
      -- 
    ca_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_1, ack => testConfigure_CP_684_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/cr
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_update_start_
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/$entry
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_609_inst_ack_0, ack => testConfigure_CP_684_elements(106)); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(106), ack => RPIPE_zeropad_input_pipe_609_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_609_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/rr
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_609_inst_ack_1, ack => testConfigure_CP_684_elements(107)); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(107), ack => type_cast_613_inst_req_0); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(107), ack => RPIPE_zeropad_input_pipe_627_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Sample/ra
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_0, ack => testConfigure_CP_684_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	131 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/ca
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_1, ack => testConfigure_CP_684_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_update_start_
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/cr
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_627_inst_ack_0, ack => testConfigure_CP_684_elements(110)); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(110), ack => RPIPE_zeropad_input_pipe_627_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_627_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/$entry
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_627_inst_ack_1, ack => testConfigure_CP_684_elements(111)); -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(111), ack => type_cast_631_inst_req_0); -- 
    rr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(111), ack => RPIPE_zeropad_input_pipe_645_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_sample_completed_
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_0, ack => testConfigure_CP_684_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	131 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_update_completed_
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_1, ack => testConfigure_CP_684_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_update_start_
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Sample/$exit
      -- 
    ra_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_645_inst_ack_0, ack => testConfigure_CP_684_elements(114)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(114), ack => RPIPE_zeropad_input_pipe_645_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_645_Update/$exit
      -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_645_inst_ack_1, ack => testConfigure_CP_684_elements(115)); -- 
    rr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(115), ack => type_cast_649_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_sample_completed_
      -- 
    ra_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => testConfigure_CP_684_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	131 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_update_completed_
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => testConfigure_CP_684_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/split_req
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/split_ack
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/$exit
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/ptr_deref_657_Split/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/rr
      -- 
    rr_1862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(118), ack => ptr_deref_657_store_0_req_0); -- 
    testConfigure_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(85) & testConfigure_CP_684_elements(89) & testConfigure_CP_684_elements(93) & testConfigure_CP_684_elements(97) & testConfigure_CP_684_elements(101) & testConfigure_CP_684_elements(105) & testConfigure_CP_684_elements(109) & testConfigure_CP_684_elements(113) & testConfigure_CP_684_elements(117);
      gj_testConfigure_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Sample/word_access_start/word_0/ra
      -- 
    ra_1863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_store_0_ack_0, ack => testConfigure_CP_684_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	131 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/$exit
      -- 
    ca_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_store_0_ack_1, ack => testConfigure_CP_684_elements(120)); -- 
    -- CP-element group 121:  branch  join  transition  place  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	82 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (10) 
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671__entry__
      -- CP-element group 121: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670__exit__
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_if_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_else_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_eval_test/branch_req
      -- CP-element group 121: 	 branch_block_stmt_277/R_exitcond7_672_place
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_dead_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_eval_test/$entry
      -- CP-element group 121: 	 branch_block_stmt_277/if_stmt_671_eval_test/$exit
      -- CP-element group 121: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/$exit
      -- 
    branch_req_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(121), ack => if_stmt_671_branch_req_0); -- 
    testConfigure_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(82) & testConfigure_CP_684_elements(120);
      gj_testConfigure_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  merge  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	132 
    -- CP-element group 122:  members (13) 
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xendx_xloopexit_forx_xend
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677__exit__
      -- CP-element group 122: 	 branch_block_stmt_277/if_stmt_671_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 122: 	 branch_block_stmt_277/if_stmt_671_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiReqMerge
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiAck/$entry
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiAck/$exit
      -- CP-element group 122: 	 branch_block_stmt_277/merge_stmt_677_PhiAck/dummy
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_277/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_671_branch_ack_1, ack => testConfigure_CP_684_elements(122)); -- 
    -- CP-element group 123:  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: 	128 
    -- CP-element group 123:  members (12) 
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody
      -- CP-element group 123: 	 branch_block_stmt_277/if_stmt_671_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/cr
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/$entry
      -- CP-element group 123: 	 branch_block_stmt_277/if_stmt_671_else_link/else_choice_transition
      -- 
    else_choice_transition_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_671_branch_ack_0, ack => testConfigure_CP_684_elements(123)); -- 
    cr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(123), ack => type_cast_514_inst_req_1); -- 
    rr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(123), ack => type_cast_514_inst_req_0); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	132 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/ra
      -- 
    ra_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_682_inst_ack_0, ack => testConfigure_CP_684_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	132 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (16) 
      -- CP-element group 125: 	 branch_block_stmt_277/branch_block_stmt_277__exit__
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685__exit__
      -- CP-element group 125: 	 branch_block_stmt_277/return__
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683__exit__
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/$exit
      -- CP-element group 125: 	 $exit
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_277/assign_stmt_683/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/return___PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_277/return___PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiReqMerge
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiAck/$entry
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiAck/$exit
      -- CP-element group 125: 	 branch_block_stmt_277/merge_stmt_685_PhiAck/dummy
      -- 
    ca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_682_inst_ack_1, ack => testConfigure_CP_684_elements(125)); -- 
    -- CP-element group 126:  transition  output  delay-element  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	81 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	130 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_req
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$exit
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_512_konst_delay_trans
      -- CP-element group 126: 	 branch_block_stmt_277/bbx_xnph_forx_xbody_PhiReq/phi_stmt_508/$exit
      -- 
    phi_stmt_508_req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_508_req_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(126), ack => phi_stmt_508_req_0); -- 
    -- Element group testConfigure_CP_684_elements(126) is a control-delay.
    cp_element_126_delay: control_delay_element  generic map(name => " 126_delay", delay_value => 1)  port map(req => testConfigure_CP_684_elements(81), ack => testConfigure_CP_684_elements(126), clk => clk, reset =>reset);
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	123 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Sample/ra
      -- 
    ra_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_514_inst_ack_0, ack => testConfigure_CP_684_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/ca
      -- CP-element group 128: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/Update/$exit
      -- 
    ca_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_514_inst_ack_1, ack => testConfigure_CP_684_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/SplitProtocol/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/type_cast_514/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_req
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/$exit
      -- CP-element group 129: 	 branch_block_stmt_277/forx_xbody_forx_xbody_PhiReq/phi_stmt_508/phi_stmt_508_sources/$exit
      -- 
    phi_stmt_508_req_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_508_req_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(129), ack => phi_stmt_508_req_1); -- 
    testConfigure_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_684_elements(127) & testConfigure_CP_684_elements(128);
      gj_testConfigure_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_684_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  transition  place  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	126 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_277/merge_stmt_507_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_277/merge_stmt_507_PhiAck/$entry
      -- 
    testConfigure_CP_684_elements(130) <= OrReduce(testConfigure_CP_684_elements(126) & testConfigure_CP_684_elements(129));
    -- CP-element group 131:  fork  transition  place  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	82 
    -- CP-element group 131: 	83 
    -- CP-element group 131: 	85 
    -- CP-element group 131: 	86 
    -- CP-element group 131: 	89 
    -- CP-element group 131: 	93 
    -- CP-element group 131: 	97 
    -- CP-element group 131: 	101 
    -- CP-element group 131: 	105 
    -- CP-element group 131: 	109 
    -- CP-element group 131: 	113 
    -- CP-element group 131: 	117 
    -- CP-element group 131: 	120 
    -- CP-element group 131:  members (56) 
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/index_resize_ack
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_update_start
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/$exit
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670__entry__
      -- CP-element group 131: 	 branch_block_stmt_277/merge_stmt_507__exit__
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/scale_rename_req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Sample/req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scale_1/scale_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_613_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_complete/req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_final_index_sum_regn_Update/req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_631_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_541_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_595_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/word_0/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_528_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/word_access_complete/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/index_resize_req
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_649_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/ptr_deref_657_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_577_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/$exit
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resize_1/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/RPIPE_zeropad_input_pipe_524_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_computed_1
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/type_cast_559_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/$entry
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/addr_of_521_update_start_
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_resized_1
      -- CP-element group 131: 	 branch_block_stmt_277/assign_stmt_522_to_assign_stmt_670/array_obj_ref_520_index_scaled_1
      -- CP-element group 131: 	 branch_block_stmt_277/merge_stmt_507_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_277/merge_stmt_507_PhiAck/phi_stmt_508_ack
      -- 
    phi_stmt_508_ack_1964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_508_ack_0, ack => testConfigure_CP_684_elements(131)); -- 
    cr_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_595_inst_req_1); -- 
    cr_1627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_528_inst_req_1); -- 
    req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => array_obj_ref_520_index_offset_req_0); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_613_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_631_inst_req_1); -- 
    req_1599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => addr_of_521_final_reg_req_1); -- 
    req_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => array_obj_ref_520_index_offset_req_1); -- 
    cr_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_541_inst_req_1); -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_649_inst_req_1); -- 
    cr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => ptr_deref_657_store_0_req_1); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_577_inst_req_1); -- 
    rr_1608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => RPIPE_zeropad_input_pipe_524_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(131), ack => type_cast_559_inst_req_1); -- 
    -- CP-element group 132:  merge  fork  transition  place  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	78 
    -- CP-element group 132: 	122 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	124 
    -- CP-element group 132: 	125 
    -- CP-element group 132:  members (13) 
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683__entry__
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679__exit__
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_update_start_
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/assign_stmt_683/type_cast_682_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiReqMerge
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiAck/$entry
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiAck/$exit
      -- CP-element group 132: 	 branch_block_stmt_277/merge_stmt_679_PhiAck/dummy
      -- 
    rr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(132), ack => type_cast_682_inst_req_0); -- 
    cr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_684_elements(132), ack => type_cast_682_inst_req_1); -- 
    testConfigure_CP_684_elements(132) <= OrReduce(testConfigure_CP_684_elements(78) & testConfigure_CP_684_elements(122));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_519_resized : std_logic_vector(13 downto 0);
    signal R_indvar_519_scaled : std_logic_vector(13 downto 0);
    signal STORE_col_high_332_data_0 : std_logic_vector(7 downto 0);
    signal STORE_col_high_332_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_depth_high_338_data_0 : std_logic_vector(7 downto 0);
    signal STORE_depth_high_338_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_pad_344_data_0 : std_logic_vector(7 downto 0);
    signal STORE_pad_344_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_row_high_326_data_0 : std_logic_vector(7 downto 0);
    signal STORE_row_high_326_word_address_0 : std_logic_vector(0 downto 0);
    signal add33_565 : std_logic_vector(63 downto 0);
    signal add39_583 : std_logic_vector(63 downto 0);
    signal add45_601 : std_logic_vector(63 downto 0);
    signal add51_619 : std_logic_vector(63 downto 0);
    signal add57_637 : std_logic_vector(63 downto 0);
    signal add63_655 : std_logic_vector(63 downto 0);
    signal add_547 : std_logic_vector(63 downto 0);
    signal array_obj_ref_520_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_520_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_522 : std_logic_vector(31 downto 0);
    signal call11_387 : std_logic_vector(7 downto 0);
    signal call1_308 : std_logic_vector(7 downto 0);
    signal call22_525 : std_logic_vector(7 downto 0);
    signal call25_538 : std_logic_vector(7 downto 0);
    signal call30_556 : std_logic_vector(7 downto 0);
    signal call36_574 : std_logic_vector(7 downto 0);
    signal call3_325 : std_logic_vector(7 downto 0);
    signal call42_592 : std_logic_vector(7 downto 0);
    signal call48_610 : std_logic_vector(7 downto 0);
    signal call4_331 : std_logic_vector(7 downto 0);
    signal call54_628 : std_logic_vector(7 downto 0);
    signal call5_337 : std_logic_vector(7 downto 0);
    signal call60_646 : std_logic_vector(7 downto 0);
    signal call6_343 : std_logic_vector(7 downto 0);
    signal call7_349 : std_logic_vector(7 downto 0);
    signal call9_368 : std_logic_vector(7 downto 0);
    signal call_291 : std_logic_vector(7 downto 0);
    signal cmp71_465 : std_logic_vector(0 downto 0);
    signal conv10_372 : std_logic_vector(31 downto 0);
    signal conv12_391 : std_logic_vector(31 downto 0);
    signal conv16_453 : std_logic_vector(63 downto 0);
    signal conv23_529 : std_logic_vector(63 downto 0);
    signal conv27_542 : std_logic_vector(63 downto 0);
    signal conv2_312 : std_logic_vector(31 downto 0);
    signal conv32_560 : std_logic_vector(63 downto 0);
    signal conv38_578 : std_logic_vector(63 downto 0);
    signal conv44_596 : std_logic_vector(63 downto 0);
    signal conv50_614 : std_logic_vector(63 downto 0);
    signal conv56_632 : std_logic_vector(63 downto 0);
    signal conv62_650 : std_logic_vector(63 downto 0);
    signal conv8_353 : std_logic_vector(31 downto 0);
    signal conv_295 : std_logic_vector(31 downto 0);
    signal exitcond7_670 : std_logic_vector(0 downto 0);
    signal iNsTr_0_283 : std_logic_vector(31 downto 0);
    signal iNsTr_17_361 : std_logic_vector(31 downto 0);
    signal iNsTr_20_380 : std_logic_vector(31 downto 0);
    signal iNsTr_23_399 : std_logic_vector(31 downto 0);
    signal iNsTr_25_411 : std_logic_vector(31 downto 0);
    signal iNsTr_26_423 : std_logic_vector(31 downto 0);
    signal iNsTr_27_435 : std_logic_vector(31 downto 0);
    signal iNsTr_3_301 : std_logic_vector(31 downto 0);
    signal iNsTr_6_318 : std_logic_vector(31 downto 0);
    signal indvar_508 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_665 : std_logic_vector(63 downto 0);
    signal mul15_449 : std_logic_vector(31 downto 0);
    signal mul_444 : std_logic_vector(31 downto 0);
    signal ptr_deref_285_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_285_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_285_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_285_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_285_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_285_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_303_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_303_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_303_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_303_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_303_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_303_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_320_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_320_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_320_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_320_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_320_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_320_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_363_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_363_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_363_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_363_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_363_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_363_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_382_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_382_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_382_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_382_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_382_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_382_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_401_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_401_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_401_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_401_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_401_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_401_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_414_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_414_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_414_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_414_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_414_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_426_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_438_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_438_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_438_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_438_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_438_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_657_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_657_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_657_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_657_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_657_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_657_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl29_553 : std_logic_vector(63 downto 0);
    signal shl35_571 : std_logic_vector(63 downto 0);
    signal shl41_589 : std_logic_vector(63 downto 0);
    signal shl47_607 : std_logic_vector(63 downto 0);
    signal shl53_625 : std_logic_vector(63 downto 0);
    signal shl59_643 : std_logic_vector(63 downto 0);
    signal shl_535 : std_logic_vector(63 downto 0);
    signal shr70x_xmask_459 : std_logic_vector(63 downto 0);
    signal tmp13_427 : std_logic_vector(31 downto 0);
    signal tmp14_439 : std_logic_vector(31 downto 0);
    signal tmp1_477 : std_logic_vector(31 downto 0);
    signal tmp2_482 : std_logic_vector(31 downto 0);
    signal tmp3_486 : std_logic_vector(63 downto 0);
    signal tmp4_492 : std_logic_vector(63 downto 0);
    signal tmp5_498 : std_logic_vector(0 downto 0);
    signal tmp_415 : std_logic_vector(31 downto 0);
    signal type_cast_287_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_490_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_503_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_514_wire : std_logic_vector(63 downto 0);
    signal type_cast_533_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_569_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_587_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_623_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_663_wire_constant : std_logic_vector(63 downto 0);
    signal umax6_505 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_col_high_332_word_address_0 <= "0";
    STORE_depth_high_338_word_address_0 <= "0";
    STORE_pad_344_word_address_0 <= "0";
    STORE_row_high_326_word_address_0 <= "0";
    array_obj_ref_520_constant_part_of_offset <= "00000000000000";
    array_obj_ref_520_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_520_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_520_resized_base_address <= "00000000000000";
    iNsTr_0_283 <= "00000000000000000000000000000000";
    iNsTr_17_361 <= "00000000000000000000000000000011";
    iNsTr_20_380 <= "00000000000000000000000000000100";
    iNsTr_23_399 <= "00000000000000000000000000000101";
    iNsTr_25_411 <= "00000000000000000000000000000011";
    iNsTr_26_423 <= "00000000000000000000000000000100";
    iNsTr_27_435 <= "00000000000000000000000000000101";
    iNsTr_3_301 <= "00000000000000000000000000000001";
    iNsTr_6_318 <= "00000000000000000000000000000010";
    ptr_deref_285_word_offset_0 <= "0000000";
    ptr_deref_303_word_offset_0 <= "0000000";
    ptr_deref_320_word_offset_0 <= "0000000";
    ptr_deref_363_word_offset_0 <= "0000000";
    ptr_deref_382_word_offset_0 <= "0000000";
    ptr_deref_401_word_offset_0 <= "0000000";
    ptr_deref_414_word_offset_0 <= "0000000";
    ptr_deref_426_word_offset_0 <= "0000000";
    ptr_deref_438_word_offset_0 <= "0000000";
    ptr_deref_657_word_offset_0 <= "00000000000000";
    type_cast_287_wire_constant <= "00000000000000000000000000000101";
    type_cast_457_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_490_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_503_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_533_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_551_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_569_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_587_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_623_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_641_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_663_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_508: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_512_wire_constant & type_cast_514_wire;
      req <= phi_stmt_508_req_0 & phi_stmt_508_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_508",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_508_ack_0,
          idata => idata,
          odata => indvar_508,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_508
    -- flow-through select operator MUX_504_inst
    umax6_505 <= tmp4_492 when (tmp5_498(0) /=  '0') else type_cast_503_wire_constant;
    addr_of_521_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_521_final_reg_req_0;
      addr_of_521_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_521_final_reg_req_1;
      addr_of_521_final_reg_ack_1<= rack(0);
      addr_of_521_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_521_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_520_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_294_inst_req_0;
      type_cast_294_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_294_inst_req_1;
      type_cast_294_inst_ack_1<= rack(0);
      type_cast_294_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_294_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_311_inst_req_0;
      type_cast_311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_311_inst_req_1;
      type_cast_311_inst_ack_1<= rack(0);
      type_cast_311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_352_inst_req_0;
      type_cast_352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_352_inst_req_1;
      type_cast_352_inst_ack_1<= rack(0);
      type_cast_352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call9_368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_390_inst_req_0;
      type_cast_390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_390_inst_req_1;
      type_cast_390_inst_ack_1<= rack(0);
      type_cast_390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul15_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_485_inst_req_0;
      type_cast_485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_485_inst_req_1;
      type_cast_485_inst_ack_1<= rack(0);
      type_cast_485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp2_482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_514_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_514_inst_req_0;
      type_cast_514_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_514_inst_req_1;
      type_cast_514_inst_ack_1<= rack(0);
      type_cast_514_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_514_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_514_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_528_inst_req_0;
      type_cast_528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_528_inst_req_1;
      type_cast_528_inst_ack_1<= rack(0);
      type_cast_528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_541_inst_req_0;
      type_cast_541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_541_inst_req_1;
      type_cast_541_inst_ack_1<= rack(0);
      type_cast_541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call25_538,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_559_inst_req_0;
      type_cast_559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_559_inst_req_1;
      type_cast_559_inst_ack_1<= rack(0);
      type_cast_559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_577_inst_req_0;
      type_cast_577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_577_inst_req_1;
      type_cast_577_inst_ack_1<= rack(0);
      type_cast_577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_595_inst_req_0;
      type_cast_595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_595_inst_req_1;
      type_cast_595_inst_ack_1<= rack(0);
      type_cast_595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_613_inst_req_0;
      type_cast_613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_613_inst_req_1;
      type_cast_613_inst_ack_1<= rack(0);
      type_cast_613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call48_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_631_inst_req_0;
      type_cast_631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_631_inst_req_1;
      type_cast_631_inst_ack_1<= rack(0);
      type_cast_631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call54_628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call60_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_682_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_682_inst_req_0;
      type_cast_682_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_682_inst_req_1;
      type_cast_682_inst_ack_1<= rack(0);
      type_cast_682_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_682_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul15_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_col_high_332_gather_scatter
    process(call4_331) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call4_331;
      ov(7 downto 0) := iv;
      STORE_col_high_332_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_depth_high_338_gather_scatter
    process(call5_337) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call5_337;
      ov(7 downto 0) := iv;
      STORE_depth_high_338_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_pad_344_gather_scatter
    process(call6_343) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call6_343;
      ov(7 downto 0) := iv;
      STORE_pad_344_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_row_high_326_gather_scatter
    process(call3_325) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call3_325;
      ov(7 downto 0) := iv;
      STORE_row_high_326_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_520_index_1_rename
    process(R_indvar_519_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_519_resized;
      ov(13 downto 0) := iv;
      R_indvar_519_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_520_index_1_resize
    process(indvar_508) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_508;
      ov := iv(13 downto 0);
      R_indvar_519_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_520_root_address_inst
    process(array_obj_ref_520_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_520_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_520_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_addr_0
    process(ptr_deref_285_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_285_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_285_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_base_resize
    process(iNsTr_0_283) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_283;
      ov := iv(6 downto 0);
      ptr_deref_285_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_gather_scatter
    process(type_cast_287_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_287_wire_constant;
      ov(31 downto 0) := iv;
      ptr_deref_285_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_285_root_address_inst
    process(ptr_deref_285_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_285_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_285_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_addr_0
    process(ptr_deref_303_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_303_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_303_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_base_resize
    process(iNsTr_3_301) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_301;
      ov := iv(6 downto 0);
      ptr_deref_303_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_gather_scatter
    process(conv_295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_295;
      ov(31 downto 0) := iv;
      ptr_deref_303_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_303_root_address_inst
    process(ptr_deref_303_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_303_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_303_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_addr_0
    process(ptr_deref_320_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_320_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_320_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_base_resize
    process(iNsTr_6_318) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_318;
      ov := iv(6 downto 0);
      ptr_deref_320_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_gather_scatter
    process(conv2_312) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv2_312;
      ov(31 downto 0) := iv;
      ptr_deref_320_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_320_root_address_inst
    process(ptr_deref_320_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_320_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_320_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_addr_0
    process(ptr_deref_363_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_363_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_363_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_base_resize
    process(iNsTr_17_361) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_17_361;
      ov := iv(6 downto 0);
      ptr_deref_363_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_gather_scatter
    process(conv8_353) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv8_353;
      ov(31 downto 0) := iv;
      ptr_deref_363_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_363_root_address_inst
    process(ptr_deref_363_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_363_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_363_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_addr_0
    process(ptr_deref_382_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_382_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_base_resize
    process(iNsTr_20_380) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_20_380;
      ov := iv(6 downto 0);
      ptr_deref_382_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_gather_scatter
    process(conv10_372) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10_372;
      ov(31 downto 0) := iv;
      ptr_deref_382_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_382_root_address_inst
    process(ptr_deref_382_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_382_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_382_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_addr_0
    process(ptr_deref_401_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_401_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_base_resize
    process(iNsTr_23_399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_23_399;
      ov := iv(6 downto 0);
      ptr_deref_401_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_gather_scatter
    process(conv12_391) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv12_391;
      ov(31 downto 0) := iv;
      ptr_deref_401_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_root_address_inst
    process(ptr_deref_401_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_401_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_addr_0
    process(ptr_deref_414_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_414_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_base_resize
    process(iNsTr_25_411) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_411;
      ov := iv(6 downto 0);
      ptr_deref_414_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_gather_scatter
    process(ptr_deref_414_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_data_0;
      ov(31 downto 0) := iv;
      tmp_415 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_414_root_address_inst
    process(ptr_deref_414_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_414_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_414_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_addr_0
    process(ptr_deref_426_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_base_resize
    process(iNsTr_26_423) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_423;
      ov := iv(6 downto 0);
      ptr_deref_426_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_gather_scatter
    process(ptr_deref_426_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_data_0;
      ov(31 downto 0) := iv;
      tmp13_427 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_root_address_inst
    process(ptr_deref_426_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_addr_0
    process(ptr_deref_438_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_438_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_base_resize
    process(iNsTr_27_435) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_27_435;
      ov := iv(6 downto 0);
      ptr_deref_438_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_gather_scatter
    process(ptr_deref_438_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_data_0;
      ov(31 downto 0) := iv;
      tmp14_439 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_438_root_address_inst
    process(ptr_deref_438_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_438_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_438_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_addr_0
    process(ptr_deref_657_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_657_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_657_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_base_resize
    process(arrayidx_522) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_522;
      ov := iv(13 downto 0);
      ptr_deref_657_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_gather_scatter
    process(add63_655) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add63_655;
      ov(63 downto 0) := iv;
      ptr_deref_657_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_657_root_address_inst
    process(ptr_deref_657_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_657_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_657_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_466_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp71_465;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_466_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_466_branch_req_0,
          ack0 => if_stmt_466_branch_ack_0,
          ack1 => if_stmt_466_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_671_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_670;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_671_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_671_branch_req_0,
          ack0 => if_stmt_671_branch_ack_0,
          ack1 => if_stmt_671_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_664_inst
    process(indvar_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_508, type_cast_663_wire_constant, tmp_var);
      indvarx_xnext_665 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_458_inst
    process(conv16_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv16_453, type_cast_457_wire_constant, tmp_var);
      shr70x_xmask_459 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_464_inst
    process(shr70x_xmask_459) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr70x_xmask_459, type_cast_463_wire_constant, tmp_var);
      cmp71_465 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_669_inst
    process(indvarx_xnext_665, umax6_505) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_665, umax6_505, tmp_var);
      exitcond7_670 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_491_inst
    process(tmp3_486) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_486, type_cast_490_wire_constant, tmp_var);
      tmp4_492 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_443_inst
    process(tmp13_427, tmp_415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_427, tmp_415, tmp_var);
      mul_444 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_448_inst
    process(mul_444, tmp14_439) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_444, tmp14_439, tmp_var);
      mul15_449 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_476_inst
    process(tmp13_427, tmp_415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_427, tmp_415, tmp_var);
      tmp1_477 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_481_inst
    process(tmp1_477, tmp14_439) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_477, tmp14_439, tmp_var);
      tmp2_482 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_546_inst
    process(shl_535, conv27_542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_535, conv27_542, tmp_var);
      add_547 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_564_inst
    process(shl29_553, conv32_560) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl29_553, conv32_560, tmp_var);
      add33_565 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_582_inst
    process(shl35_571, conv38_578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl35_571, conv38_578, tmp_var);
      add39_583 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_600_inst
    process(shl41_589, conv44_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl41_589, conv44_596, tmp_var);
      add45_601 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_618_inst
    process(shl47_607, conv50_614) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl47_607, conv50_614, tmp_var);
      add51_619 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_636_inst
    process(shl53_625, conv56_632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl53_625, conv56_632, tmp_var);
      add57_637 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_654_inst
    process(shl59_643, conv62_650) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl59_643, conv62_650, tmp_var);
      add63_655 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_534_inst
    process(conv23_529) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv23_529, type_cast_533_wire_constant, tmp_var);
      shl_535 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_552_inst
    process(add_547) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_547, type_cast_551_wire_constant, tmp_var);
      shl29_553 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_570_inst
    process(add33_565) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add33_565, type_cast_569_wire_constant, tmp_var);
      shl35_571 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_588_inst
    process(add39_583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add39_583, type_cast_587_wire_constant, tmp_var);
      shl41_589 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_606_inst
    process(add45_601) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add45_601, type_cast_605_wire_constant, tmp_var);
      shl47_607 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_624_inst
    process(add51_619) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add51_619, type_cast_623_wire_constant, tmp_var);
      shl53_625 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_642_inst
    process(add57_637) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_637, type_cast_641_wire_constant, tmp_var);
      shl59_643 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_497_inst
    process(tmp4_492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp4_492, type_cast_496_wire_constant, tmp_var);
      tmp5_498 <= tmp_var; --
    end process;
    -- shared split operator group (24) : array_obj_ref_520_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_519_scaled;
      array_obj_ref_520_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_520_index_offset_req_0;
      array_obj_ref_520_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_520_index_offset_req_1;
      array_obj_ref_520_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_414_load_0 ptr_deref_426_load_0 ptr_deref_438_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_414_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_426_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_438_load_0_req_0;
      ptr_deref_414_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_426_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_438_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_414_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_426_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_438_load_0_req_1;
      ptr_deref_414_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_426_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_438_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_414_word_address_0 & ptr_deref_426_word_address_0 & ptr_deref_438_word_address_0;
      ptr_deref_414_data_0 <= data_out(95 downto 64);
      ptr_deref_426_data_0 <= data_out(63 downto 32);
      ptr_deref_438_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(6 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : STORE_col_high_332_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_col_high_332_store_0_req_0;
      STORE_col_high_332_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_col_high_332_store_0_req_1;
      STORE_col_high_332_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_col_high_332_word_address_0;
      data_in <= STORE_col_high_332_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_depth_high_338_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_depth_high_338_store_0_req_0;
      STORE_depth_high_338_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_depth_high_338_store_0_req_1;
      STORE_depth_high_338_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_depth_high_338_word_address_0;
      data_in <= STORE_depth_high_338_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_pad_344_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_pad_344_store_0_req_0;
      STORE_pad_344_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_pad_344_store_0_req_1;
      STORE_pad_344_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_pad_344_word_address_0;
      data_in <= STORE_pad_344_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : STORE_row_high_326_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_row_high_326_store_0_req_0;
      STORE_row_high_326_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_row_high_326_store_0_req_1;
      STORE_row_high_326_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_row_high_326_word_address_0;
      data_in <= STORE_row_high_326_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_285_store_0 ptr_deref_303_store_0 ptr_deref_320_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_285_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_303_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_320_store_0_req_0;
      ptr_deref_285_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_303_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_320_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_285_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_303_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_320_store_0_req_1;
      ptr_deref_285_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_303_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_320_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_285_word_address_0 & ptr_deref_303_word_address_0 & ptr_deref_320_word_address_0;
      data_in <= ptr_deref_285_data_0 & ptr_deref_303_data_0 & ptr_deref_320_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(6 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_363_store_0 ptr_deref_382_store_0 ptr_deref_401_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_363_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_382_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_401_store_0_req_0;
      ptr_deref_363_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_382_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_401_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_363_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_382_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_401_store_0_req_1;
      ptr_deref_363_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_382_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_401_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_363_word_address_0 & ptr_deref_382_word_address_0 & ptr_deref_401_word_address_0;
      data_in <= ptr_deref_363_data_0 & ptr_deref_382_data_0 & ptr_deref_401_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(6 downto 0),
          mdata => memory_space_6_sr_data(31 downto 0),
          mtag => memory_space_6_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_657_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_657_store_0_req_0;
      ptr_deref_657_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_657_store_0_req_1;
      ptr_deref_657_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_657_word_address_0;
      data_in <= ptr_deref_657_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_627_inst RPIPE_zeropad_input_pipe_645_inst RPIPE_zeropad_input_pipe_609_inst RPIPE_zeropad_input_pipe_591_inst RPIPE_zeropad_input_pipe_573_inst RPIPE_zeropad_input_pipe_290_inst RPIPE_zeropad_input_pipe_307_inst RPIPE_zeropad_input_pipe_324_inst RPIPE_zeropad_input_pipe_330_inst RPIPE_zeropad_input_pipe_336_inst RPIPE_zeropad_input_pipe_342_inst RPIPE_zeropad_input_pipe_348_inst RPIPE_zeropad_input_pipe_367_inst RPIPE_zeropad_input_pipe_386_inst RPIPE_zeropad_input_pipe_524_inst RPIPE_zeropad_input_pipe_537_inst RPIPE_zeropad_input_pipe_555_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(135 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 16 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_627_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_645_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_609_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_591_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_573_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_290_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_307_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_324_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_330_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_336_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_342_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_348_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_367_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_386_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_524_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_537_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_555_inst_req_0;
      RPIPE_zeropad_input_pipe_627_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_645_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_609_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_591_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_573_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_290_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_307_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_324_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_330_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_336_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_342_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_348_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_367_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_386_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_524_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_537_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_555_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_627_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_645_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_609_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_591_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_573_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_290_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_307_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_324_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_330_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_336_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_342_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_348_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_367_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_386_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_524_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_537_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_555_inst_req_1;
      RPIPE_zeropad_input_pipe_627_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_645_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_609_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_591_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_573_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_290_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_307_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_324_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_330_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_336_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_342_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_348_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_367_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_386_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_524_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_537_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_555_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      call54_628 <= data_out(135 downto 128);
      call60_646 <= data_out(127 downto 120);
      call48_610 <= data_out(119 downto 112);
      call42_592 <= data_out(111 downto 104);
      call36_574 <= data_out(103 downto 96);
      call_291 <= data_out(95 downto 88);
      call1_308 <= data_out(87 downto 80);
      call3_325 <= data_out(79 downto 72);
      call4_331 <= data_out(71 downto 64);
      call5_337 <= data_out(63 downto 56);
      call6_343 <= data_out(55 downto 48);
      call7_349 <= data_out(47 downto 40);
      call9_368 <= data_out(39 downto 32);
      call11_387 <= data_out(31 downto 24);
      call22_525 <= data_out(23 downto 16);
      call25_538 <= data_out(15 downto 8);
      call30_556 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 17,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_2152_start: Boolean;
  signal zeropad3D_CP_2152_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ptr_deref_1076_store_0_req_1 : boolean;
  signal if_stmt_984_branch_req_0 : boolean;
  signal type_cast_1031_inst_req_0 : boolean;
  signal LOAD_row_high_941_load_0_ack_0 : boolean;
  signal type_cast_975_inst_ack_1 : boolean;
  signal type_cast_975_inst_req_1 : boolean;
  signal type_cast_1031_inst_ack_0 : boolean;
  signal if_stmt_984_branch_ack_1 : boolean;
  signal type_cast_1149_inst_req_1 : boolean;
  signal type_cast_1149_inst_ack_1 : boolean;
  signal call_stmt_716_call_req_0 : boolean;
  signal call_stmt_716_call_ack_0 : boolean;
  signal call_stmt_716_call_req_1 : boolean;
  signal call_stmt_716_call_ack_1 : boolean;
  signal ptr_deref_727_load_0_req_0 : boolean;
  signal ptr_deref_727_load_0_ack_0 : boolean;
  signal ptr_deref_727_load_0_req_1 : boolean;
  signal ptr_deref_727_load_0_ack_1 : boolean;
  signal type_cast_731_inst_req_0 : boolean;
  signal type_cast_731_inst_ack_0 : boolean;
  signal type_cast_731_inst_req_1 : boolean;
  signal type_cast_731_inst_ack_1 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal STORE_row_high_733_store_0_req_0 : boolean;
  signal STORE_row_high_733_store_0_ack_0 : boolean;
  signal STORE_row_high_733_store_0_req_1 : boolean;
  signal if_stmt_1016_branch_ack_0 : boolean;
  signal STORE_row_high_733_store_0_ack_1 : boolean;
  signal array_obj_ref_1711_index_offset_ack_0 : boolean;
  signal if_stmt_1016_branch_ack_1 : boolean;
  signal type_cast_975_inst_ack_0 : boolean;
  signal type_cast_975_inst_req_0 : boolean;
  signal ptr_deref_746_load_0_req_0 : boolean;
  signal ptr_deref_746_load_0_ack_0 : boolean;
  signal LOAD_row_high_941_load_0_req_0 : boolean;
  signal ptr_deref_746_load_0_req_1 : boolean;
  signal ptr_deref_746_load_0_ack_1 : boolean;
  signal type_cast_1149_inst_ack_0 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal if_stmt_1016_branch_req_0 : boolean;
  signal type_cast_1149_inst_req_0 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal ptr_deref_1160_load_0_ack_1 : boolean;
  signal STORE_col_high_752_store_0_req_0 : boolean;
  signal STORE_col_high_752_store_0_ack_0 : boolean;
  signal STORE_col_high_752_store_0_req_1 : boolean;
  signal STORE_col_high_752_store_0_ack_1 : boolean;
  signal type_cast_1174_inst_ack_1 : boolean;
  signal LOAD_row_high_941_load_0_ack_1 : boolean;
  signal type_cast_996_inst_ack_1 : boolean;
  signal type_cast_996_inst_req_1 : boolean;
  signal ptr_deref_765_load_0_req_0 : boolean;
  signal ptr_deref_765_load_0_ack_0 : boolean;
  signal if_stmt_965_branch_ack_0 : boolean;
  signal ptr_deref_765_load_0_req_1 : boolean;
  signal type_cast_996_inst_ack_0 : boolean;
  signal ptr_deref_765_load_0_ack_1 : boolean;
  signal type_cast_996_inst_req_0 : boolean;
  signal addr_of_1156_final_reg_ack_1 : boolean;
  signal addr_of_1156_final_reg_req_1 : boolean;
  signal type_cast_769_inst_req_0 : boolean;
  signal type_cast_769_inst_ack_0 : boolean;
  signal type_cast_1085_inst_ack_1 : boolean;
  signal type_cast_769_inst_req_1 : boolean;
  signal type_cast_1066_inst_ack_1 : boolean;
  signal type_cast_769_inst_ack_1 : boolean;
  signal ptr_deref_1160_load_0_req_1 : boolean;
  signal addr_of_1156_final_reg_ack_0 : boolean;
  signal addr_of_1156_final_reg_req_0 : boolean;
  signal type_cast_1085_inst_req_1 : boolean;
  signal type_cast_1066_inst_req_1 : boolean;
  signal STORE_depth_high_771_store_0_req_0 : boolean;
  signal STORE_depth_high_771_store_0_ack_0 : boolean;
  signal LOAD_row_high_941_load_0_req_1 : boolean;
  signal STORE_depth_high_771_store_0_req_1 : boolean;
  signal STORE_depth_high_771_store_0_ack_1 : boolean;
  signal type_cast_1174_inst_req_1 : boolean;
  signal ptr_deref_1076_store_0_ack_0 : boolean;
  signal ptr_deref_1076_store_0_req_0 : boolean;
  signal addr_of_1073_final_reg_ack_1 : boolean;
  signal type_cast_1026_inst_ack_1 : boolean;
  signal addr_of_1073_final_reg_req_1 : boolean;
  signal if_stmt_965_branch_ack_1 : boolean;
  signal LOAD_pad_776_load_0_req_0 : boolean;
  signal LOAD_pad_776_load_0_ack_0 : boolean;
  signal type_cast_1026_inst_req_1 : boolean;
  signal LOAD_pad_776_load_0_req_1 : boolean;
  signal LOAD_pad_776_load_0_ack_1 : boolean;
  signal LOAD_col_high_992_load_0_ack_1 : boolean;
  signal type_cast_1085_inst_ack_0 : boolean;
  signal LOAD_depth_high_779_load_0_req_0 : boolean;
  signal LOAD_col_high_992_load_0_req_1 : boolean;
  signal LOAD_depth_high_779_load_0_ack_0 : boolean;
  signal if_stmt_965_branch_req_0 : boolean;
  signal LOAD_depth_high_779_load_0_req_1 : boolean;
  signal LOAD_depth_high_779_load_0_ack_1 : boolean;
  signal type_cast_1085_inst_req_0 : boolean;
  signal LOAD_col_high_782_load_0_req_0 : boolean;
  signal LOAD_col_high_992_load_0_ack_0 : boolean;
  signal LOAD_col_high_782_load_0_ack_0 : boolean;
  signal LOAD_col_high_992_load_0_req_0 : boolean;
  signal LOAD_col_high_782_load_0_req_1 : boolean;
  signal LOAD_col_high_782_load_0_ack_1 : boolean;
  signal addr_of_1073_final_reg_ack_0 : boolean;
  signal addr_of_1073_final_reg_req_0 : boolean;
  signal type_cast_1066_inst_ack_0 : boolean;
  signal type_cast_1066_inst_req_0 : boolean;
  signal ptr_deref_1160_load_0_ack_0 : boolean;
  signal ptr_deref_794_load_0_req_0 : boolean;
  signal ptr_deref_794_load_0_ack_0 : boolean;
  signal type_cast_1026_inst_ack_0 : boolean;
  signal type_cast_945_inst_ack_1 : boolean;
  signal ptr_deref_794_load_0_req_1 : boolean;
  signal ptr_deref_794_load_0_ack_1 : boolean;
  signal type_cast_945_inst_req_1 : boolean;
  signal array_obj_ref_1155_index_offset_ack_1 : boolean;
  signal array_obj_ref_1155_index_offset_req_1 : boolean;
  signal array_obj_ref_1072_index_offset_ack_1 : boolean;
  signal array_obj_ref_1072_index_offset_req_1 : boolean;
  signal array_obj_ref_1072_index_offset_ack_0 : boolean;
  signal array_obj_ref_1072_index_offset_req_0 : boolean;
  signal ptr_deref_1160_load_0_req_0 : boolean;
  signal type_cast_1026_inst_req_0 : boolean;
  signal type_cast_945_inst_ack_0 : boolean;
  signal ptr_deref_806_load_0_req_0 : boolean;
  signal ptr_deref_806_load_0_ack_0 : boolean;
  signal type_cast_945_inst_req_0 : boolean;
  signal ptr_deref_806_load_0_req_1 : boolean;
  signal ptr_deref_806_load_0_ack_1 : boolean;
  signal type_cast_810_inst_req_0 : boolean;
  signal type_cast_810_inst_ack_0 : boolean;
  signal if_stmt_933_branch_ack_0 : boolean;
  signal type_cast_810_inst_req_1 : boolean;
  signal type_cast_1031_inst_ack_1 : boolean;
  signal type_cast_810_inst_ack_1 : boolean;
  signal array_obj_ref_1155_index_offset_ack_0 : boolean;
  signal array_obj_ref_1155_index_offset_req_0 : boolean;
  signal if_stmt_984_branch_ack_0 : boolean;
  signal type_cast_1031_inst_req_1 : boolean;
  signal type_cast_814_inst_req_0 : boolean;
  signal type_cast_814_inst_ack_0 : boolean;
  signal ptr_deref_1076_store_0_ack_1 : boolean;
  signal type_cast_814_inst_req_1 : boolean;
  signal type_cast_814_inst_ack_1 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal array_obj_ref_1628_index_offset_req_1 : boolean;
  signal type_cast_924_inst_req_0 : boolean;
  signal array_obj_ref_1628_index_offset_ack_1 : boolean;
  signal type_cast_924_inst_ack_0 : boolean;
  signal type_cast_924_inst_req_1 : boolean;
  signal type_cast_924_inst_ack_1 : boolean;
  signal if_stmt_933_branch_req_0 : boolean;
  signal if_stmt_933_branch_ack_1 : boolean;
  signal array_obj_ref_1180_index_offset_req_0 : boolean;
  signal array_obj_ref_1180_index_offset_ack_0 : boolean;
  signal array_obj_ref_1180_index_offset_req_1 : boolean;
  signal array_obj_ref_1180_index_offset_ack_1 : boolean;
  signal addr_of_1181_final_reg_req_0 : boolean;
  signal addr_of_1181_final_reg_ack_0 : boolean;
  signal addr_of_1181_final_reg_req_1 : boolean;
  signal addr_of_1181_final_reg_ack_1 : boolean;
  signal type_cast_1641_inst_ack_0 : boolean;
  signal type_cast_1641_inst_req_0 : boolean;
  signal LOAD_col_high_1555_load_0_ack_1 : boolean;
  signal ptr_deref_1184_store_0_req_0 : boolean;
  signal ptr_deref_1184_store_0_ack_0 : boolean;
  signal LOAD_col_high_1555_load_0_req_1 : boolean;
  signal ptr_deref_1184_store_0_req_1 : boolean;
  signal ptr_deref_1184_store_0_ack_1 : boolean;
  signal addr_of_1737_final_reg_req_1 : boolean;
  signal array_obj_ref_2269_index_offset_req_1 : boolean;
  signal type_cast_1559_inst_ack_0 : boolean;
  signal array_obj_ref_1628_index_offset_ack_0 : boolean;
  signal array_obj_ref_1711_index_offset_req_0 : boolean;
  signal type_cast_1192_inst_req_0 : boolean;
  signal type_cast_1192_inst_ack_0 : boolean;
  signal type_cast_1192_inst_req_1 : boolean;
  signal type_cast_1192_inst_ack_1 : boolean;
  signal array_obj_ref_1628_index_offset_req_0 : boolean;
  signal ptr_deref_1716_load_0_ack_0 : boolean;
  signal ptr_deref_1716_load_0_req_0 : boolean;
  signal if_stmt_1207_branch_req_0 : boolean;
  signal if_stmt_1207_branch_ack_1 : boolean;
  signal if_stmt_1207_branch_ack_0 : boolean;
  signal addr_of_1712_final_reg_ack_0 : boolean;
  signal addr_of_1712_final_reg_req_0 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal array_obj_ref_1736_index_offset_ack_0 : boolean;
  signal LOAD_col_high_1555_load_0_ack_0 : boolean;
  signal LOAD_col_high_1555_load_0_req_0 : boolean;
  signal LOAD_col_high_1234_load_0_req_0 : boolean;
  signal LOAD_col_high_1234_load_0_ack_0 : boolean;
  signal LOAD_col_high_1234_load_0_req_1 : boolean;
  signal LOAD_col_high_1234_load_0_ack_1 : boolean;
  signal ptr_deref_1632_store_0_ack_1 : boolean;
  signal ptr_deref_1632_store_0_req_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal array_obj_ref_1736_index_offset_req_0 : boolean;
  signal addr_of_1737_final_reg_ack_0 : boolean;
  signal type_cast_1258_inst_req_0 : boolean;
  signal type_cast_1258_inst_ack_0 : boolean;
  signal type_cast_1258_inst_req_1 : boolean;
  signal type_cast_1258_inst_ack_1 : boolean;
  signal addr_of_1737_final_reg_req_0 : boolean;
  signal type_cast_1275_inst_req_0 : boolean;
  signal ptr_deref_1632_store_0_ack_0 : boolean;
  signal type_cast_1275_inst_ack_0 : boolean;
  signal addr_of_1629_final_reg_ack_1 : boolean;
  signal type_cast_1275_inst_req_1 : boolean;
  signal ptr_deref_1632_store_0_req_0 : boolean;
  signal type_cast_1275_inst_ack_1 : boolean;
  signal type_cast_1730_inst_ack_1 : boolean;
  signal LOAD_row_high_1278_load_0_req_0 : boolean;
  signal LOAD_row_high_1278_load_0_ack_0 : boolean;
  signal LOAD_row_high_1278_load_0_req_1 : boolean;
  signal LOAD_row_high_1278_load_0_ack_1 : boolean;
  signal addr_of_1629_final_reg_req_1 : boolean;
  signal if_stmt_1547_branch_ack_0 : boolean;
  signal type_cast_1282_inst_req_0 : boolean;
  signal type_cast_1282_inst_ack_0 : boolean;
  signal type_cast_1282_inst_req_1 : boolean;
  signal type_cast_1282_inst_ack_1 : boolean;
  signal type_cast_1730_inst_req_1 : boolean;
  signal array_obj_ref_1736_index_offset_ack_1 : boolean;
  signal if_stmt_1300_branch_req_0 : boolean;
  signal if_stmt_1300_branch_ack_1 : boolean;
  signal if_stmt_1300_branch_ack_0 : boolean;
  signal addr_of_1629_final_reg_ack_0 : boolean;
  signal addr_of_1629_final_reg_req_0 : boolean;
  signal if_stmt_1573_branch_ack_0 : boolean;
  signal LOAD_col_high_1331_load_0_req_0 : boolean;
  signal LOAD_col_high_1331_load_0_ack_0 : boolean;
  signal LOAD_col_high_1331_load_0_req_1 : boolean;
  signal type_cast_1622_inst_ack_1 : boolean;
  signal LOAD_col_high_1331_load_0_ack_1 : boolean;
  signal type_cast_1622_inst_req_1 : boolean;
  signal ptr_deref_1716_load_0_ack_1 : boolean;
  signal array_obj_ref_1736_index_offset_req_1 : boolean;
  signal ptr_deref_1716_load_0_req_1 : boolean;
  signal array_obj_ref_1711_index_offset_ack_1 : boolean;
  signal type_cast_1335_inst_req_0 : boolean;
  signal type_cast_1335_inst_ack_0 : boolean;
  signal type_cast_1335_inst_req_1 : boolean;
  signal type_cast_1335_inst_ack_1 : boolean;
  signal type_cast_1730_inst_ack_0 : boolean;
  signal LOAD_pad_1344_load_0_req_0 : boolean;
  signal type_cast_1622_inst_ack_0 : boolean;
  signal LOAD_pad_1344_load_0_ack_0 : boolean;
  signal if_stmt_1573_branch_ack_1 : boolean;
  signal LOAD_pad_1344_load_0_req_1 : boolean;
  signal type_cast_1622_inst_req_0 : boolean;
  signal LOAD_pad_1344_load_0_ack_1 : boolean;
  signal type_cast_1730_inst_req_0 : boolean;
  signal array_obj_ref_1711_index_offset_req_1 : boolean;
  signal LOAD_depth_high_1347_load_0_req_0 : boolean;
  signal LOAD_depth_high_1347_load_0_ack_0 : boolean;
  signal LOAD_depth_high_1347_load_0_req_1 : boolean;
  signal type_cast_1588_inst_ack_1 : boolean;
  signal LOAD_depth_high_1347_load_0_ack_1 : boolean;
  signal type_cast_1588_inst_req_1 : boolean;
  signal type_cast_1705_inst_ack_1 : boolean;
  signal type_cast_1705_inst_req_1 : boolean;
  signal type_cast_1588_inst_ack_0 : boolean;
  signal if_stmt_1573_branch_req_0 : boolean;
  signal ptr_deref_1359_load_0_req_0 : boolean;
  signal type_cast_1588_inst_req_0 : boolean;
  signal ptr_deref_1359_load_0_ack_0 : boolean;
  signal ptr_deref_1359_load_0_req_1 : boolean;
  signal ptr_deref_1359_load_0_ack_1 : boolean;
  signal addr_of_1737_final_reg_ack_1 : boolean;
  signal type_cast_1705_inst_ack_0 : boolean;
  signal type_cast_1705_inst_req_0 : boolean;
  signal type_cast_1559_inst_ack_1 : boolean;
  signal ptr_deref_1371_load_0_req_0 : boolean;
  signal type_cast_1583_inst_ack_1 : boolean;
  signal ptr_deref_1371_load_0_ack_0 : boolean;
  signal if_stmt_1547_branch_ack_1 : boolean;
  signal type_cast_1559_inst_req_1 : boolean;
  signal ptr_deref_1371_load_0_req_1 : boolean;
  signal type_cast_1583_inst_req_1 : boolean;
  signal ptr_deref_1371_load_0_ack_1 : boolean;
  signal type_cast_1559_inst_req_0 : boolean;
  signal type_cast_1583_inst_ack_0 : boolean;
  signal type_cast_1583_inst_req_0 : boolean;
  signal type_cast_1375_inst_req_0 : boolean;
  signal type_cast_1375_inst_ack_0 : boolean;
  signal addr_of_1712_final_reg_ack_1 : boolean;
  signal type_cast_1375_inst_req_1 : boolean;
  signal type_cast_1375_inst_ack_1 : boolean;
  signal type_cast_1641_inst_ack_1 : boolean;
  signal type_cast_1641_inst_req_1 : boolean;
  signal type_cast_1379_inst_req_0 : boolean;
  signal type_cast_1379_inst_ack_0 : boolean;
  signal addr_of_1712_final_reg_req_1 : boolean;
  signal type_cast_1379_inst_req_1 : boolean;
  signal type_cast_1379_inst_ack_1 : boolean;
  signal array_obj_ref_2269_index_offset_ack_1 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal type_cast_2141_inst_req_0 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_2146_inst_req_1 : boolean;
  signal type_cast_1487_inst_req_0 : boolean;
  signal type_cast_1487_inst_ack_0 : boolean;
  signal type_cast_1487_inst_req_1 : boolean;
  signal type_cast_1487_inst_ack_1 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal type_cast_2146_inst_ack_1 : boolean;
  signal type_cast_2180_inst_ack_0 : boolean;
  signal if_stmt_1496_branch_req_0 : boolean;
  signal if_stmt_1496_branch_ack_1 : boolean;
  signal type_cast_2141_inst_ack_0 : boolean;
  signal if_stmt_1496_branch_ack_0 : boolean;
  signal LOAD_row_high_1504_load_0_req_0 : boolean;
  signal LOAD_row_high_1504_load_0_ack_0 : boolean;
  signal LOAD_row_high_1504_load_0_req_1 : boolean;
  signal LOAD_row_high_1504_load_0_ack_1 : boolean;
  signal type_cast_1508_inst_req_0 : boolean;
  signal type_cast_1508_inst_ack_0 : boolean;
  signal type_cast_1508_inst_req_1 : boolean;
  signal type_cast_1508_inst_ack_1 : boolean;
  signal if_stmt_1528_branch_req_0 : boolean;
  signal if_stmt_1528_branch_ack_1 : boolean;
  signal if_stmt_1528_branch_ack_0 : boolean;
  signal type_cast_1538_inst_req_0 : boolean;
  signal type_cast_1538_inst_ack_0 : boolean;
  signal type_cast_1538_inst_req_1 : boolean;
  signal type_cast_1538_inst_ack_1 : boolean;
  signal if_stmt_1547_branch_req_0 : boolean;
  signal phi_stmt_4704_req_1 : boolean;
  signal phi_stmt_4145_ack_0 : boolean;
  signal ptr_deref_1740_store_0_req_0 : boolean;
  signal ptr_deref_1740_store_0_ack_0 : boolean;
  signal ptr_deref_1740_store_0_req_1 : boolean;
  signal ptr_deref_1740_store_0_ack_1 : boolean;
  signal type_cast_1748_inst_req_0 : boolean;
  signal type_cast_1748_inst_ack_0 : boolean;
  signal type_cast_1748_inst_req_1 : boolean;
  signal type_cast_1748_inst_ack_1 : boolean;
  signal if_stmt_1763_branch_req_0 : boolean;
  signal if_stmt_1763_branch_ack_1 : boolean;
  signal if_stmt_1763_branch_ack_0 : boolean;
  signal type_cast_1787_inst_req_0 : boolean;
  signal type_cast_1787_inst_ack_0 : boolean;
  signal type_cast_1787_inst_req_1 : boolean;
  signal type_cast_1787_inst_ack_1 : boolean;
  signal addr_of_2295_final_reg_ack_1 : boolean;
  signal addr_of_2295_final_reg_ack_0 : boolean;
  signal addr_of_2295_final_reg_req_0 : boolean;
  signal ptr_deref_2274_load_0_ack_0 : boolean;
  signal ptr_deref_2190_store_0_ack_0 : boolean;
  signal ptr_deref_2190_store_0_req_0 : boolean;
  signal LOAD_col_high_1790_load_0_req_0 : boolean;
  signal LOAD_col_high_1790_load_0_ack_0 : boolean;
  signal LOAD_col_high_1790_load_0_req_1 : boolean;
  signal LOAD_col_high_1790_load_0_ack_1 : boolean;
  signal type_cast_1794_inst_req_0 : boolean;
  signal array_obj_ref_2269_index_offset_ack_0 : boolean;
  signal type_cast_1794_inst_ack_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_1794_inst_req_1 : boolean;
  signal array_obj_ref_2269_index_offset_req_0 : boolean;
  signal type_cast_1794_inst_ack_1 : boolean;
  signal addr_of_2295_final_reg_req_1 : boolean;
  signal type_cast_2288_inst_ack_1 : boolean;
  signal type_cast_1808_inst_req_0 : boolean;
  signal type_cast_1808_inst_ack_0 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2288_inst_req_1 : boolean;
  signal type_cast_1808_inst_req_1 : boolean;
  signal type_cast_1808_inst_ack_1 : boolean;
  signal type_cast_1824_inst_req_0 : boolean;
  signal type_cast_1824_inst_ack_0 : boolean;
  signal type_cast_2288_inst_ack_0 : boolean;
  signal type_cast_1824_inst_req_1 : boolean;
  signal type_cast_1824_inst_ack_1 : boolean;
  signal type_cast_2146_inst_ack_0 : boolean;
  signal type_cast_2146_inst_req_0 : boolean;
  signal LOAD_row_high_1827_load_0_req_0 : boolean;
  signal LOAD_row_high_1827_load_0_ack_0 : boolean;
  signal LOAD_row_high_1827_load_0_req_1 : boolean;
  signal LOAD_row_high_1827_load_0_ack_1 : boolean;
  signal type_cast_2288_inst_req_0 : boolean;
  signal type_cast_1831_inst_req_0 : boolean;
  signal type_cast_1831_inst_ack_0 : boolean;
  signal type_cast_1831_inst_req_1 : boolean;
  signal type_cast_1831_inst_ack_1 : boolean;
  signal array_obj_ref_2294_index_offset_ack_1 : boolean;
  signal array_obj_ref_2294_index_offset_req_1 : boolean;
  signal if_stmt_1849_branch_req_0 : boolean;
  signal if_stmt_1849_branch_ack_1 : boolean;
  signal if_stmt_1849_branch_ack_0 : boolean;
  signal ptr_deref_2274_load_0_req_0 : boolean;
  signal LOAD_row_high_1880_load_0_req_0 : boolean;
  signal LOAD_row_high_1880_load_0_ack_0 : boolean;
  signal LOAD_row_high_1880_load_0_req_1 : boolean;
  signal LOAD_row_high_1880_load_0_ack_1 : boolean;
  signal type_cast_1884_inst_req_0 : boolean;
  signal type_cast_1884_inst_ack_0 : boolean;
  signal ptr_deref_2190_store_0_ack_1 : boolean;
  signal type_cast_1884_inst_req_1 : boolean;
  signal type_cast_1884_inst_ack_1 : boolean;
  signal type_cast_2141_inst_ack_1 : boolean;
  signal LOAD_pad_1893_load_0_req_0 : boolean;
  signal LOAD_pad_1893_load_0_ack_0 : boolean;
  signal type_cast_2141_inst_req_1 : boolean;
  signal LOAD_pad_1893_load_0_req_1 : boolean;
  signal LOAD_pad_1893_load_0_ack_1 : boolean;
  signal array_obj_ref_2294_index_offset_ack_0 : boolean;
  signal array_obj_ref_2294_index_offset_req_0 : boolean;
  signal ptr_deref_2274_load_0_ack_1 : boolean;
  signal LOAD_depth_high_1896_load_0_req_0 : boolean;
  signal LOAD_depth_high_1896_load_0_ack_0 : boolean;
  signal LOAD_depth_high_1896_load_0_req_1 : boolean;
  signal LOAD_depth_high_1896_load_0_ack_1 : boolean;
  signal ptr_deref_2190_store_0_req_1 : boolean;
  signal ptr_deref_2274_load_0_req_1 : boolean;
  signal LOAD_col_high_1899_load_0_req_0 : boolean;
  signal LOAD_col_high_1899_load_0_ack_0 : boolean;
  signal LOAD_col_high_1899_load_0_req_1 : boolean;
  signal addr_of_2187_final_reg_ack_1 : boolean;
  signal LOAD_col_high_1899_load_0_ack_1 : boolean;
  signal addr_of_2187_final_reg_req_1 : boolean;
  signal addr_of_2270_final_reg_ack_1 : boolean;
  signal addr_of_2270_final_reg_req_1 : boolean;
  signal addr_of_2270_final_reg_ack_0 : boolean;
  signal type_cast_2263_inst_ack_1 : boolean;
  signal type_cast_2263_inst_req_1 : boolean;
  signal addr_of_2187_final_reg_ack_0 : boolean;
  signal addr_of_2187_final_reg_req_0 : boolean;
  signal ptr_deref_1911_load_0_req_0 : boolean;
  signal ptr_deref_1911_load_0_ack_0 : boolean;
  signal ptr_deref_1911_load_0_req_1 : boolean;
  signal ptr_deref_1911_load_0_ack_1 : boolean;
  signal type_cast_2180_inst_req_0 : boolean;
  signal addr_of_2270_final_reg_req_0 : boolean;
  signal array_obj_ref_2186_index_offset_ack_1 : boolean;
  signal array_obj_ref_2186_index_offset_req_1 : boolean;
  signal type_cast_2263_inst_ack_0 : boolean;
  signal array_obj_ref_2186_index_offset_ack_0 : boolean;
  signal type_cast_2263_inst_req_0 : boolean;
  signal array_obj_ref_2186_index_offset_req_0 : boolean;
  signal if_stmt_2131_branch_ack_0 : boolean;
  signal type_cast_2180_inst_ack_1 : boolean;
  signal type_cast_2180_inst_req_1 : boolean;
  signal ptr_deref_1923_load_0_req_0 : boolean;
  signal ptr_deref_1923_load_0_ack_0 : boolean;
  signal ptr_deref_1923_load_0_req_1 : boolean;
  signal ptr_deref_1923_load_0_ack_1 : boolean;
  signal type_cast_1927_inst_req_0 : boolean;
  signal type_cast_1927_inst_ack_0 : boolean;
  signal type_cast_1927_inst_req_1 : boolean;
  signal type_cast_1927_inst_ack_1 : boolean;
  signal type_cast_1931_inst_req_0 : boolean;
  signal type_cast_1931_inst_ack_0 : boolean;
  signal type_cast_1931_inst_req_1 : boolean;
  signal type_cast_1931_inst_ack_1 : boolean;
  signal type_cast_1970_inst_req_0 : boolean;
  signal type_cast_1970_inst_ack_0 : boolean;
  signal type_cast_1970_inst_req_1 : boolean;
  signal type_cast_1970_inst_ack_1 : boolean;
  signal type_cast_2039_inst_req_0 : boolean;
  signal type_cast_2039_inst_ack_0 : boolean;
  signal type_cast_2039_inst_req_1 : boolean;
  signal type_cast_2039_inst_ack_1 : boolean;
  signal if_stmt_2048_branch_req_0 : boolean;
  signal if_stmt_2048_branch_ack_1 : boolean;
  signal if_stmt_2048_branch_ack_0 : boolean;
  signal LOAD_row_high_2056_load_0_req_0 : boolean;
  signal addr_of_2838_final_reg_req_0 : boolean;
  signal LOAD_row_high_2056_load_0_ack_0 : boolean;
  signal LOAD_row_high_2056_load_0_req_1 : boolean;
  signal LOAD_row_high_2056_load_0_ack_1 : boolean;
  signal addr_of_2838_final_reg_ack_0 : boolean;
  signal addr_of_2755_final_reg_req_0 : boolean;
  signal type_cast_2060_inst_req_0 : boolean;
  signal type_cast_2060_inst_ack_0 : boolean;
  signal type_cast_2060_inst_req_1 : boolean;
  signal type_cast_2060_inst_ack_1 : boolean;
  signal if_stmt_2080_branch_req_0 : boolean;
  signal if_stmt_2080_branch_ack_1 : boolean;
  signal if_stmt_2080_branch_ack_0 : boolean;
  signal type_cast_2090_inst_req_0 : boolean;
  signal type_cast_2090_inst_ack_0 : boolean;
  signal type_cast_2090_inst_req_1 : boolean;
  signal type_cast_2090_inst_ack_1 : boolean;
  signal if_stmt_2099_branch_req_0 : boolean;
  signal if_stmt_2099_branch_ack_1 : boolean;
  signal if_stmt_2099_branch_ack_0 : boolean;
  signal LOAD_col_high_2107_load_0_req_0 : boolean;
  signal LOAD_col_high_2107_load_0_ack_0 : boolean;
  signal LOAD_col_high_2107_load_0_req_1 : boolean;
  signal LOAD_col_high_2107_load_0_ack_1 : boolean;
  signal type_cast_2111_inst_req_0 : boolean;
  signal type_cast_2111_inst_ack_0 : boolean;
  signal type_cast_2111_inst_req_1 : boolean;
  signal type_cast_2111_inst_ack_1 : boolean;
  signal if_stmt_2131_branch_req_0 : boolean;
  signal if_stmt_2131_branch_ack_1 : boolean;
  signal ptr_deref_2298_store_0_req_0 : boolean;
  signal ptr_deref_2298_store_0_ack_0 : boolean;
  signal ptr_deref_2298_store_0_req_1 : boolean;
  signal ptr_deref_2298_store_0_ack_1 : boolean;
  signal type_cast_2306_inst_req_0 : boolean;
  signal type_cast_2306_inst_ack_0 : boolean;
  signal type_cast_2306_inst_req_1 : boolean;
  signal type_cast_2306_inst_ack_1 : boolean;
  signal if_stmt_2321_branch_req_0 : boolean;
  signal if_stmt_2321_branch_ack_1 : boolean;
  signal if_stmt_2321_branch_ack_0 : boolean;
  signal type_cast_2345_inst_req_0 : boolean;
  signal type_cast_2345_inst_ack_0 : boolean;
  signal type_cast_2345_inst_req_1 : boolean;
  signal type_cast_2345_inst_ack_1 : boolean;
  signal LOAD_col_high_2348_load_0_req_0 : boolean;
  signal LOAD_col_high_2348_load_0_ack_0 : boolean;
  signal LOAD_col_high_2348_load_0_req_1 : boolean;
  signal LOAD_col_high_2348_load_0_ack_1 : boolean;
  signal type_cast_2352_inst_req_0 : boolean;
  signal type_cast_2352_inst_ack_0 : boolean;
  signal type_cast_2352_inst_req_1 : boolean;
  signal type_cast_2352_inst_ack_1 : boolean;
  signal array_obj_ref_2862_index_offset_ack_0 : boolean;
  signal type_cast_2372_inst_req_0 : boolean;
  signal ptr_deref_2842_load_0_ack_1 : boolean;
  signal type_cast_2372_inst_ack_0 : boolean;
  signal array_obj_ref_2862_index_offset_req_0 : boolean;
  signal type_cast_2372_inst_req_1 : boolean;
  signal ptr_deref_2842_load_0_req_1 : boolean;
  signal type_cast_2372_inst_ack_1 : boolean;
  signal addr_of_2863_final_reg_ack_1 : boolean;
  signal type_cast_2856_inst_ack_1 : boolean;
  signal type_cast_2389_inst_req_0 : boolean;
  signal type_cast_2389_inst_ack_0 : boolean;
  signal type_cast_2389_inst_req_1 : boolean;
  signal type_cast_2389_inst_ack_1 : boolean;
  signal addr_of_2863_final_reg_req_1 : boolean;
  signal type_cast_2856_inst_req_1 : boolean;
  signal array_obj_ref_2837_index_offset_ack_1 : boolean;
  signal array_obj_ref_2837_index_offset_req_1 : boolean;
  signal array_obj_ref_2837_index_offset_ack_0 : boolean;
  signal LOAD_row_high_2392_load_0_req_0 : boolean;
  signal array_obj_ref_2837_index_offset_req_0 : boolean;
  signal LOAD_row_high_2392_load_0_ack_0 : boolean;
  signal LOAD_row_high_2392_load_0_req_1 : boolean;
  signal LOAD_row_high_2392_load_0_ack_1 : boolean;
  signal addr_of_2863_final_reg_ack_0 : boolean;
  signal type_cast_2396_inst_req_0 : boolean;
  signal type_cast_2396_inst_ack_0 : boolean;
  signal type_cast_2396_inst_req_1 : boolean;
  signal type_cast_2396_inst_ack_1 : boolean;
  signal array_obj_ref_2754_index_offset_ack_1 : boolean;
  signal array_obj_ref_2754_index_offset_req_1 : boolean;
  signal ptr_deref_2842_load_0_ack_0 : boolean;
  signal if_stmt_2414_branch_req_0 : boolean;
  signal ptr_deref_2842_load_0_req_0 : boolean;
  signal if_stmt_2414_branch_ack_1 : boolean;
  signal if_stmt_2414_branch_ack_0 : boolean;
  signal array_obj_ref_2754_index_offset_ack_0 : boolean;
  signal addr_of_2838_final_reg_ack_1 : boolean;
  signal LOAD_col_high_2445_load_0_req_0 : boolean;
  signal LOAD_col_high_2445_load_0_ack_0 : boolean;
  signal LOAD_col_high_2445_load_0_req_1 : boolean;
  signal LOAD_col_high_2445_load_0_ack_1 : boolean;
  signal addr_of_2838_final_reg_req_1 : boolean;
  signal addr_of_2863_final_reg_req_0 : boolean;
  signal type_cast_2449_inst_req_0 : boolean;
  signal type_cast_2449_inst_ack_0 : boolean;
  signal type_cast_2449_inst_req_1 : boolean;
  signal type_cast_2449_inst_ack_1 : boolean;
  signal type_cast_2856_inst_ack_0 : boolean;
  signal type_cast_2856_inst_req_0 : boolean;
  signal LOAD_row_high_2458_load_0_req_0 : boolean;
  signal LOAD_row_high_2458_load_0_ack_0 : boolean;
  signal LOAD_row_high_2458_load_0_req_1 : boolean;
  signal LOAD_row_high_2458_load_0_ack_1 : boolean;
  signal type_cast_2831_inst_ack_1 : boolean;
  signal type_cast_2831_inst_req_1 : boolean;
  signal type_cast_2831_inst_ack_0 : boolean;
  signal type_cast_2831_inst_req_0 : boolean;
  signal type_cast_2462_inst_req_0 : boolean;
  signal type_cast_2462_inst_ack_0 : boolean;
  signal type_cast_2462_inst_req_1 : boolean;
  signal type_cast_2462_inst_ack_1 : boolean;
  signal type_cast_3395_inst_ack_1 : boolean;
  signal array_obj_ref_2754_index_offset_req_0 : boolean;
  signal LOAD_pad_2471_load_0_req_0 : boolean;
  signal LOAD_pad_2471_load_0_ack_0 : boolean;
  signal LOAD_pad_2471_load_0_req_1 : boolean;
  signal LOAD_pad_2471_load_0_ack_1 : boolean;
  signal type_cast_2767_inst_ack_1 : boolean;
  signal type_cast_2767_inst_req_1 : boolean;
  signal LOAD_depth_high_2474_load_0_req_0 : boolean;
  signal type_cast_2767_inst_ack_0 : boolean;
  signal LOAD_depth_high_2474_load_0_ack_0 : boolean;
  signal type_cast_2767_inst_req_0 : boolean;
  signal LOAD_depth_high_2474_load_0_req_1 : boolean;
  signal LOAD_depth_high_2474_load_0_ack_1 : boolean;
  signal array_obj_ref_2862_index_offset_ack_1 : boolean;
  signal array_obj_ref_2862_index_offset_req_1 : boolean;
  signal ptr_deref_2758_store_0_ack_1 : boolean;
  signal ptr_deref_2758_store_0_req_1 : boolean;
  signal addr_of_2755_final_reg_ack_1 : boolean;
  signal addr_of_2755_final_reg_req_1 : boolean;
  signal ptr_deref_2758_store_0_ack_0 : boolean;
  signal ptr_deref_2486_load_0_req_0 : boolean;
  signal ptr_deref_2758_store_0_req_0 : boolean;
  signal ptr_deref_2486_load_0_ack_0 : boolean;
  signal ptr_deref_2486_load_0_req_1 : boolean;
  signal ptr_deref_2486_load_0_ack_1 : boolean;
  signal array_obj_ref_3426_index_offset_req_1 : boolean;
  signal addr_of_2755_final_reg_ack_0 : boolean;
  signal array_obj_ref_3426_index_offset_req_0 : boolean;
  signal array_obj_ref_3426_index_offset_ack_1 : boolean;
  signal ptr_deref_2498_load_0_req_0 : boolean;
  signal ptr_deref_2498_load_0_ack_0 : boolean;
  signal ptr_deref_2498_load_0_req_1 : boolean;
  signal ptr_deref_2498_load_0_ack_1 : boolean;
  signal addr_of_3427_final_reg_ack_1 : boolean;
  signal ptr_deref_3322_store_0_req_0 : boolean;
  signal type_cast_2502_inst_req_0 : boolean;
  signal ptr_deref_3406_load_0_req_1 : boolean;
  signal type_cast_2502_inst_ack_0 : boolean;
  signal ptr_deref_3322_store_0_ack_0 : boolean;
  signal type_cast_2502_inst_req_1 : boolean;
  signal type_cast_2502_inst_ack_1 : boolean;
  signal ptr_deref_3406_load_0_ack_1 : boolean;
  signal type_cast_2506_inst_req_0 : boolean;
  signal type_cast_2506_inst_ack_0 : boolean;
  signal type_cast_2506_inst_req_1 : boolean;
  signal type_cast_2506_inst_ack_1 : boolean;
  signal type_cast_2545_inst_req_0 : boolean;
  signal type_cast_2545_inst_ack_0 : boolean;
  signal type_cast_2545_inst_req_1 : boolean;
  signal type_cast_2545_inst_ack_1 : boolean;
  signal type_cast_2613_inst_req_0 : boolean;
  signal type_cast_2613_inst_ack_0 : boolean;
  signal type_cast_3420_inst_req_0 : boolean;
  signal type_cast_2613_inst_req_1 : boolean;
  signal type_cast_2613_inst_ack_1 : boolean;
  signal type_cast_3331_inst_req_1 : boolean;
  signal if_stmt_2622_branch_req_0 : boolean;
  signal type_cast_3331_inst_ack_1 : boolean;
  signal if_stmt_2622_branch_ack_1 : boolean;
  signal if_stmt_2622_branch_ack_0 : boolean;
  signal type_cast_3420_inst_ack_0 : boolean;
  signal array_obj_ref_3426_index_offset_ack_0 : boolean;
  signal LOAD_row_high_2630_load_0_req_0 : boolean;
  signal LOAD_row_high_2630_load_0_ack_0 : boolean;
  signal LOAD_row_high_2630_load_0_req_1 : boolean;
  signal LOAD_row_high_2630_load_0_ack_1 : boolean;
  signal ptr_deref_3322_store_0_req_1 : boolean;
  signal type_cast_2634_inst_req_0 : boolean;
  signal type_cast_2634_inst_ack_0 : boolean;
  signal ptr_deref_3322_store_0_ack_1 : boolean;
  signal type_cast_2634_inst_req_1 : boolean;
  signal type_cast_2634_inst_ack_1 : boolean;
  signal if_stmt_2654_branch_req_0 : boolean;
  signal if_stmt_2654_branch_ack_1 : boolean;
  signal if_stmt_2654_branch_ack_0 : boolean;
  signal type_cast_3420_inst_req_1 : boolean;
  signal type_cast_2664_inst_req_0 : boolean;
  signal type_cast_2664_inst_ack_0 : boolean;
  signal type_cast_2664_inst_req_1 : boolean;
  signal type_cast_2664_inst_ack_1 : boolean;
  signal if_stmt_2673_branch_req_0 : boolean;
  signal if_stmt_2673_branch_ack_1 : boolean;
  signal if_stmt_2673_branch_ack_0 : boolean;
  signal LOAD_col_high_2681_load_0_req_0 : boolean;
  signal LOAD_col_high_2681_load_0_ack_0 : boolean;
  signal LOAD_col_high_2681_load_0_req_1 : boolean;
  signal LOAD_col_high_2681_load_0_ack_1 : boolean;
  signal type_cast_2685_inst_req_0 : boolean;
  signal type_cast_2685_inst_ack_0 : boolean;
  signal type_cast_2685_inst_req_1 : boolean;
  signal type_cast_2685_inst_ack_1 : boolean;
  signal if_stmt_2699_branch_req_0 : boolean;
  signal if_stmt_2699_branch_ack_1 : boolean;
  signal if_stmt_2699_branch_ack_0 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal type_cast_2714_inst_req_0 : boolean;
  signal type_cast_2714_inst_ack_0 : boolean;
  signal type_cast_2714_inst_req_1 : boolean;
  signal type_cast_2714_inst_ack_1 : boolean;
  signal type_cast_2748_inst_req_0 : boolean;
  signal type_cast_2748_inst_ack_0 : boolean;
  signal type_cast_2748_inst_req_1 : boolean;
  signal type_cast_2748_inst_ack_1 : boolean;
  signal ptr_deref_2866_store_0_req_0 : boolean;
  signal ptr_deref_2866_store_0_ack_0 : boolean;
  signal ptr_deref_2866_store_0_req_1 : boolean;
  signal ptr_deref_2866_store_0_ack_1 : boolean;
  signal type_cast_2874_inst_req_0 : boolean;
  signal type_cast_2874_inst_ack_0 : boolean;
  signal type_cast_2874_inst_req_1 : boolean;
  signal type_cast_2874_inst_ack_1 : boolean;
  signal if_stmt_2889_branch_req_0 : boolean;
  signal if_stmt_2889_branch_ack_1 : boolean;
  signal if_stmt_2889_branch_ack_0 : boolean;
  signal type_cast_2913_inst_req_0 : boolean;
  signal type_cast_2913_inst_ack_0 : boolean;
  signal type_cast_2913_inst_req_1 : boolean;
  signal type_cast_2913_inst_ack_1 : boolean;
  signal LOAD_col_high_2916_load_0_req_0 : boolean;
  signal LOAD_col_high_2916_load_0_ack_0 : boolean;
  signal LOAD_col_high_2916_load_0_req_1 : boolean;
  signal LOAD_col_high_2916_load_0_ack_1 : boolean;
  signal type_cast_2920_inst_req_0 : boolean;
  signal type_cast_2920_inst_ack_0 : boolean;
  signal type_cast_2920_inst_req_1 : boolean;
  signal type_cast_2920_inst_ack_1 : boolean;
  signal type_cast_2934_inst_req_0 : boolean;
  signal type_cast_2934_inst_ack_0 : boolean;
  signal type_cast_2934_inst_req_1 : boolean;
  signal type_cast_2934_inst_ack_1 : boolean;
  signal type_cast_2950_inst_req_0 : boolean;
  signal type_cast_2950_inst_ack_0 : boolean;
  signal type_cast_2950_inst_req_1 : boolean;
  signal type_cast_2950_inst_ack_1 : boolean;
  signal LOAD_row_high_2953_load_0_req_0 : boolean;
  signal LOAD_row_high_2953_load_0_ack_0 : boolean;
  signal LOAD_row_high_2953_load_0_req_1 : boolean;
  signal LOAD_row_high_2953_load_0_ack_1 : boolean;
  signal ptr_deref_3406_load_0_ack_0 : boolean;
  signal ptr_deref_3406_load_0_req_0 : boolean;
  signal addr_of_3427_final_reg_req_1 : boolean;
  signal type_cast_2957_inst_req_0 : boolean;
  signal type_cast_2957_inst_ack_0 : boolean;
  signal type_cast_2957_inst_req_1 : boolean;
  signal type_cast_2957_inst_ack_1 : boolean;
  signal type_cast_3395_inst_req_1 : boolean;
  signal addr_of_3427_final_reg_ack_0 : boolean;
  signal if_stmt_2975_branch_req_0 : boolean;
  signal if_stmt_2975_branch_ack_1 : boolean;
  signal if_stmt_2975_branch_ack_0 : boolean;
  signal addr_of_4007_final_reg_ack_1 : boolean;
  signal type_cast_3331_inst_ack_0 : boolean;
  signal type_cast_3331_inst_req_0 : boolean;
  signal LOAD_row_high_3006_load_0_req_0 : boolean;
  signal LOAD_row_high_3006_load_0_ack_0 : boolean;
  signal LOAD_row_high_3006_load_0_req_1 : boolean;
  signal LOAD_row_high_3006_load_0_ack_1 : boolean;
  signal addr_of_3427_final_reg_req_0 : boolean;
  signal type_cast_3010_inst_req_0 : boolean;
  signal type_cast_3010_inst_ack_0 : boolean;
  signal type_cast_3010_inst_req_1 : boolean;
  signal type_cast_3010_inst_ack_1 : boolean;
  signal type_cast_3395_inst_ack_0 : boolean;
  signal type_cast_3395_inst_req_0 : boolean;
  signal LOAD_pad_3019_load_0_req_0 : boolean;
  signal LOAD_pad_3019_load_0_ack_0 : boolean;
  signal LOAD_pad_3019_load_0_req_1 : boolean;
  signal LOAD_pad_3019_load_0_ack_1 : boolean;
  signal LOAD_depth_high_3022_load_0_req_0 : boolean;
  signal LOAD_depth_high_3022_load_0_ack_0 : boolean;
  signal LOAD_depth_high_3022_load_0_req_1 : boolean;
  signal LOAD_depth_high_3022_load_0_ack_1 : boolean;
  signal addr_of_3402_final_reg_ack_1 : boolean;
  signal addr_of_3402_final_reg_req_1 : boolean;
  signal addr_of_3402_final_reg_ack_0 : boolean;
  signal addr_of_3402_final_reg_req_0 : boolean;
  signal LOAD_col_high_3025_load_0_req_0 : boolean;
  signal LOAD_col_high_3025_load_0_ack_0 : boolean;
  signal LOAD_col_high_3025_load_0_req_1 : boolean;
  signal LOAD_col_high_3025_load_0_ack_1 : boolean;
  signal array_obj_ref_3401_index_offset_ack_1 : boolean;
  signal array_obj_ref_3401_index_offset_req_1 : boolean;
  signal array_obj_ref_3401_index_offset_ack_0 : boolean;
  signal array_obj_ref_3401_index_offset_req_0 : boolean;
  signal type_cast_3420_inst_ack_1 : boolean;
  signal ptr_deref_3037_load_0_req_0 : boolean;
  signal ptr_deref_3037_load_0_ack_0 : boolean;
  signal ptr_deref_3037_load_0_req_1 : boolean;
  signal ptr_deref_3037_load_0_ack_1 : boolean;
  signal ptr_deref_3986_load_0_req_1 : boolean;
  signal addr_of_4007_final_reg_req_0 : boolean;
  signal ptr_deref_3986_load_0_ack_1 : boolean;
  signal addr_of_4007_final_reg_ack_0 : boolean;
  signal type_cast_4000_inst_req_1 : boolean;
  signal ptr_deref_3049_load_0_req_0 : boolean;
  signal ptr_deref_3049_load_0_ack_0 : boolean;
  signal ptr_deref_3049_load_0_req_1 : boolean;
  signal ptr_deref_3049_load_0_ack_1 : boolean;
  signal type_cast_3053_inst_req_0 : boolean;
  signal type_cast_3053_inst_ack_0 : boolean;
  signal type_cast_3053_inst_req_1 : boolean;
  signal type_cast_3053_inst_ack_1 : boolean;
  signal type_cast_3057_inst_req_0 : boolean;
  signal type_cast_3057_inst_ack_0 : boolean;
  signal type_cast_3057_inst_req_1 : boolean;
  signal type_cast_3057_inst_ack_1 : boolean;
  signal type_cast_4000_inst_ack_1 : boolean;
  signal array_obj_ref_4006_index_offset_req_0 : boolean;
  signal type_cast_3096_inst_req_0 : boolean;
  signal array_obj_ref_4006_index_offset_ack_0 : boolean;
  signal type_cast_3096_inst_ack_0 : boolean;
  signal type_cast_3096_inst_req_1 : boolean;
  signal type_cast_3096_inst_ack_1 : boolean;
  signal addr_of_3982_final_reg_req_1 : boolean;
  signal type_cast_3165_inst_req_0 : boolean;
  signal type_cast_3165_inst_ack_0 : boolean;
  signal type_cast_3165_inst_req_1 : boolean;
  signal type_cast_3165_inst_ack_1 : boolean;
  signal addr_of_3982_final_reg_ack_1 : boolean;
  signal if_stmt_3174_branch_req_0 : boolean;
  signal if_stmt_3174_branch_ack_1 : boolean;
  signal if_stmt_3174_branch_ack_0 : boolean;
  signal LOAD_row_high_3182_load_0_req_0 : boolean;
  signal LOAD_row_high_3182_load_0_ack_0 : boolean;
  signal LOAD_row_high_3182_load_0_req_1 : boolean;
  signal LOAD_row_high_3182_load_0_ack_1 : boolean;
  signal type_cast_4000_inst_req_0 : boolean;
  signal type_cast_4000_inst_ack_0 : boolean;
  signal type_cast_3186_inst_req_0 : boolean;
  signal array_obj_ref_4006_index_offset_req_1 : boolean;
  signal type_cast_3186_inst_ack_0 : boolean;
  signal type_cast_3186_inst_req_1 : boolean;
  signal type_cast_3186_inst_ack_1 : boolean;
  signal if_stmt_3212_branch_req_0 : boolean;
  signal if_stmt_3212_branch_ack_1 : boolean;
  signal if_stmt_3212_branch_ack_0 : boolean;
  signal type_cast_3222_inst_req_0 : boolean;
  signal array_obj_ref_4006_index_offset_ack_1 : boolean;
  signal type_cast_3222_inst_ack_0 : boolean;
  signal type_cast_3222_inst_req_1 : boolean;
  signal type_cast_3222_inst_ack_1 : boolean;
  signal if_stmt_3231_branch_req_0 : boolean;
  signal if_stmt_3231_branch_ack_1 : boolean;
  signal if_stmt_3231_branch_ack_0 : boolean;
  signal LOAD_col_high_3239_load_0_req_0 : boolean;
  signal LOAD_col_high_3239_load_0_ack_0 : boolean;
  signal LOAD_col_high_3239_load_0_req_1 : boolean;
  signal LOAD_col_high_3239_load_0_ack_1 : boolean;
  signal type_cast_3243_inst_req_0 : boolean;
  signal type_cast_3243_inst_ack_0 : boolean;
  signal type_cast_3243_inst_req_1 : boolean;
  signal type_cast_3243_inst_ack_1 : boolean;
  signal if_stmt_3263_branch_req_0 : boolean;
  signal if_stmt_3263_branch_ack_1 : boolean;
  signal if_stmt_3263_branch_ack_0 : boolean;
  signal type_cast_3273_inst_req_0 : boolean;
  signal type_cast_3273_inst_ack_0 : boolean;
  signal type_cast_3273_inst_req_1 : boolean;
  signal type_cast_3273_inst_ack_1 : boolean;
  signal type_cast_3278_inst_req_0 : boolean;
  signal type_cast_3278_inst_ack_0 : boolean;
  signal type_cast_3278_inst_req_1 : boolean;
  signal type_cast_3278_inst_ack_1 : boolean;
  signal type_cast_3312_inst_req_0 : boolean;
  signal type_cast_3312_inst_ack_0 : boolean;
  signal type_cast_3312_inst_req_1 : boolean;
  signal type_cast_3312_inst_ack_1 : boolean;
  signal array_obj_ref_3318_index_offset_req_0 : boolean;
  signal array_obj_ref_3318_index_offset_ack_0 : boolean;
  signal array_obj_ref_3318_index_offset_req_1 : boolean;
  signal array_obj_ref_3318_index_offset_ack_1 : boolean;
  signal addr_of_3319_final_reg_req_0 : boolean;
  signal addr_of_3319_final_reg_ack_0 : boolean;
  signal addr_of_3319_final_reg_req_1 : boolean;
  signal addr_of_3319_final_reg_ack_1 : boolean;
  signal ptr_deref_3430_store_0_req_0 : boolean;
  signal ptr_deref_3430_store_0_ack_0 : boolean;
  signal ptr_deref_3430_store_0_req_1 : boolean;
  signal ptr_deref_3430_store_0_ack_1 : boolean;
  signal type_cast_3438_inst_req_0 : boolean;
  signal type_cast_3438_inst_ack_0 : boolean;
  signal type_cast_3438_inst_req_1 : boolean;
  signal type_cast_3438_inst_ack_1 : boolean;
  signal if_stmt_3453_branch_req_0 : boolean;
  signal if_stmt_3453_branch_ack_1 : boolean;
  signal if_stmt_3453_branch_ack_0 : boolean;
  signal type_cast_3477_inst_req_0 : boolean;
  signal type_cast_3477_inst_ack_0 : boolean;
  signal type_cast_3477_inst_req_1 : boolean;
  signal type_cast_3477_inst_ack_1 : boolean;
  signal LOAD_col_high_3480_load_0_req_0 : boolean;
  signal LOAD_col_high_3480_load_0_ack_0 : boolean;
  signal LOAD_col_high_3480_load_0_req_1 : boolean;
  signal LOAD_col_high_3480_load_0_ack_1 : boolean;
  signal type_cast_3484_inst_req_0 : boolean;
  signal type_cast_3484_inst_ack_0 : boolean;
  signal type_cast_3484_inst_req_1 : boolean;
  signal type_cast_3484_inst_ack_1 : boolean;
  signal type_cast_3504_inst_req_0 : boolean;
  signal type_cast_3504_inst_ack_0 : boolean;
  signal type_cast_3504_inst_req_1 : boolean;
  signal type_cast_3504_inst_ack_1 : boolean;
  signal type_cast_3521_inst_req_0 : boolean;
  signal type_cast_3521_inst_ack_0 : boolean;
  signal type_cast_3521_inst_req_1 : boolean;
  signal type_cast_3521_inst_ack_1 : boolean;
  signal LOAD_row_high_3524_load_0_req_0 : boolean;
  signal LOAD_row_high_3524_load_0_ack_0 : boolean;
  signal LOAD_row_high_3524_load_0_req_1 : boolean;
  signal LOAD_row_high_3524_load_0_ack_1 : boolean;
  signal type_cast_3528_inst_req_0 : boolean;
  signal type_cast_3528_inst_ack_0 : boolean;
  signal type_cast_3528_inst_req_1 : boolean;
  signal type_cast_3528_inst_ack_1 : boolean;
  signal if_stmt_3552_branch_req_0 : boolean;
  signal if_stmt_3552_branch_ack_1 : boolean;
  signal if_stmt_3552_branch_ack_0 : boolean;
  signal LOAD_col_high_3583_load_0_req_0 : boolean;
  signal LOAD_col_high_3583_load_0_ack_0 : boolean;
  signal LOAD_col_high_3583_load_0_req_1 : boolean;
  signal LOAD_col_high_3583_load_0_ack_1 : boolean;
  signal addr_of_4007_final_reg_req_1 : boolean;
  signal ptr_deref_3986_load_0_ack_0 : boolean;
  signal type_cast_3587_inst_req_0 : boolean;
  signal type_cast_3587_inst_ack_0 : boolean;
  signal type_cast_3587_inst_req_1 : boolean;
  signal type_cast_3587_inst_ack_1 : boolean;
  signal array_obj_ref_3981_index_offset_ack_1 : boolean;
  signal array_obj_ref_3981_index_offset_req_1 : boolean;
  signal array_obj_ref_3981_index_offset_ack_0 : boolean;
  signal array_obj_ref_3981_index_offset_req_0 : boolean;
  signal LOAD_row_high_3596_load_0_req_0 : boolean;
  signal LOAD_row_high_3596_load_0_ack_0 : boolean;
  signal LOAD_row_high_3596_load_0_req_1 : boolean;
  signal LOAD_row_high_3596_load_0_ack_1 : boolean;
  signal ptr_deref_3986_load_0_req_0 : boolean;
  signal type_cast_3600_inst_req_0 : boolean;
  signal type_cast_3600_inst_ack_0 : boolean;
  signal type_cast_3600_inst_req_1 : boolean;
  signal type_cast_3600_inst_ack_1 : boolean;
  signal addr_of_3982_final_reg_ack_0 : boolean;
  signal LOAD_pad_3609_load_0_req_0 : boolean;
  signal LOAD_pad_3609_load_0_ack_0 : boolean;
  signal LOAD_pad_3609_load_0_req_1 : boolean;
  signal LOAD_pad_3609_load_0_ack_1 : boolean;
  signal addr_of_3982_final_reg_req_0 : boolean;
  signal LOAD_depth_high_3612_load_0_req_0 : boolean;
  signal LOAD_depth_high_3612_load_0_ack_0 : boolean;
  signal LOAD_depth_high_3612_load_0_req_1 : boolean;
  signal LOAD_depth_high_3612_load_0_ack_1 : boolean;
  signal addr_of_4571_final_reg_req_0 : boolean;
  signal type_cast_4564_inst_req_0 : boolean;
  signal type_cast_4564_inst_ack_0 : boolean;
  signal ptr_deref_3624_load_0_req_0 : boolean;
  signal ptr_deref_3624_load_0_ack_0 : boolean;
  signal ptr_deref_4574_store_0_req_1 : boolean;
  signal ptr_deref_3624_load_0_req_1 : boolean;
  signal ptr_deref_3624_load_0_ack_1 : boolean;
  signal addr_of_4571_final_reg_ack_0 : boolean;
  signal addr_of_4571_final_reg_req_1 : boolean;
  signal type_cast_4564_inst_req_1 : boolean;
  signal ptr_deref_3636_load_0_req_0 : boolean;
  signal ptr_deref_3636_load_0_ack_0 : boolean;
  signal type_cast_4564_inst_ack_1 : boolean;
  signal array_obj_ref_4570_index_offset_req_1 : boolean;
  signal ptr_deref_3636_load_0_req_1 : boolean;
  signal ptr_deref_3636_load_0_ack_1 : boolean;
  signal ptr_deref_4574_store_0_ack_1 : boolean;
  signal array_obj_ref_4570_index_offset_ack_1 : boolean;
  signal type_cast_3640_inst_req_0 : boolean;
  signal type_cast_3640_inst_ack_0 : boolean;
  signal type_cast_3640_inst_req_1 : boolean;
  signal type_cast_3640_inst_ack_1 : boolean;
  signal addr_of_4571_final_reg_ack_1 : boolean;
  signal type_cast_3644_inst_req_0 : boolean;
  signal type_cast_3644_inst_ack_0 : boolean;
  signal type_cast_3644_inst_req_1 : boolean;
  signal type_cast_3644_inst_ack_1 : boolean;
  signal type_cast_3683_inst_req_0 : boolean;
  signal type_cast_3683_inst_ack_0 : boolean;
  signal type_cast_3683_inst_req_1 : boolean;
  signal type_cast_3683_inst_ack_1 : boolean;
  signal type_cast_4582_inst_req_0 : boolean;
  signal type_cast_3751_inst_req_0 : boolean;
  signal type_cast_3751_inst_ack_0 : boolean;
  signal type_cast_3751_inst_req_1 : boolean;
  signal type_cast_3751_inst_ack_1 : boolean;
  signal ptr_deref_4550_load_0_req_0 : boolean;
  signal ptr_deref_4550_load_0_ack_0 : boolean;
  signal ptr_deref_4574_store_0_req_0 : boolean;
  signal if_stmt_3760_branch_req_0 : boolean;
  signal if_stmt_3760_branch_ack_1 : boolean;
  signal if_stmt_3760_branch_ack_0 : boolean;
  signal ptr_deref_4574_store_0_ack_0 : boolean;
  signal LOAD_row_high_3768_load_0_req_0 : boolean;
  signal LOAD_row_high_3768_load_0_ack_0 : boolean;
  signal LOAD_row_high_3768_load_0_req_1 : boolean;
  signal LOAD_row_high_3768_load_0_ack_1 : boolean;
  signal type_cast_3772_inst_req_0 : boolean;
  signal type_cast_3772_inst_ack_0 : boolean;
  signal type_cast_3772_inst_req_1 : boolean;
  signal type_cast_3772_inst_ack_1 : boolean;
  signal array_obj_ref_4570_index_offset_req_0 : boolean;
  signal if_stmt_3798_branch_req_0 : boolean;
  signal if_stmt_3798_branch_ack_1 : boolean;
  signal if_stmt_3798_branch_ack_0 : boolean;
  signal type_cast_3808_inst_req_0 : boolean;
  signal type_cast_3808_inst_ack_0 : boolean;
  signal type_cast_3808_inst_req_1 : boolean;
  signal type_cast_3808_inst_ack_1 : boolean;
  signal array_obj_ref_4570_index_offset_ack_0 : boolean;
  signal type_cast_4582_inst_ack_0 : boolean;
  signal if_stmt_3817_branch_req_0 : boolean;
  signal if_stmt_3817_branch_ack_1 : boolean;
  signal if_stmt_3817_branch_ack_0 : boolean;
  signal LOAD_col_high_3825_load_0_req_0 : boolean;
  signal LOAD_col_high_3825_load_0_ack_0 : boolean;
  signal LOAD_col_high_3825_load_0_req_1 : boolean;
  signal LOAD_col_high_3825_load_0_ack_1 : boolean;
  signal type_cast_3829_inst_req_0 : boolean;
  signal type_cast_3829_inst_ack_0 : boolean;
  signal type_cast_3829_inst_req_1 : boolean;
  signal type_cast_3829_inst_ack_1 : boolean;
  signal if_stmt_3843_branch_req_0 : boolean;
  signal if_stmt_3843_branch_ack_1 : boolean;
  signal if_stmt_3843_branch_ack_0 : boolean;
  signal type_cast_3853_inst_req_0 : boolean;
  signal type_cast_3853_inst_ack_0 : boolean;
  signal type_cast_3853_inst_req_1 : boolean;
  signal type_cast_3853_inst_ack_1 : boolean;
  signal type_cast_3858_inst_req_0 : boolean;
  signal type_cast_3858_inst_ack_0 : boolean;
  signal type_cast_3858_inst_req_1 : boolean;
  signal type_cast_3858_inst_ack_1 : boolean;
  signal type_cast_3892_inst_req_0 : boolean;
  signal type_cast_3892_inst_ack_0 : boolean;
  signal type_cast_3892_inst_req_1 : boolean;
  signal type_cast_3892_inst_ack_1 : boolean;
  signal array_obj_ref_3898_index_offset_req_0 : boolean;
  signal array_obj_ref_3898_index_offset_ack_0 : boolean;
  signal array_obj_ref_3898_index_offset_req_1 : boolean;
  signal array_obj_ref_3898_index_offset_ack_1 : boolean;
  signal addr_of_3899_final_reg_req_0 : boolean;
  signal addr_of_3899_final_reg_ack_0 : boolean;
  signal addr_of_3899_final_reg_req_1 : boolean;
  signal addr_of_3899_final_reg_ack_1 : boolean;
  signal ptr_deref_3902_store_0_req_0 : boolean;
  signal ptr_deref_3902_store_0_ack_0 : boolean;
  signal ptr_deref_3902_store_0_req_1 : boolean;
  signal ptr_deref_3902_store_0_ack_1 : boolean;
  signal type_cast_3911_inst_req_0 : boolean;
  signal type_cast_3911_inst_ack_0 : boolean;
  signal type_cast_3911_inst_req_1 : boolean;
  signal type_cast_3911_inst_ack_1 : boolean;
  signal type_cast_3975_inst_req_0 : boolean;
  signal type_cast_3975_inst_ack_0 : boolean;
  signal type_cast_3975_inst_req_1 : boolean;
  signal type_cast_3975_inst_ack_1 : boolean;
  signal ptr_deref_4010_store_0_req_0 : boolean;
  signal ptr_deref_4010_store_0_ack_0 : boolean;
  signal ptr_deref_4010_store_0_req_1 : boolean;
  signal ptr_deref_4010_store_0_ack_1 : boolean;
  signal type_cast_4018_inst_req_0 : boolean;
  signal type_cast_4018_inst_ack_0 : boolean;
  signal type_cast_4018_inst_req_1 : boolean;
  signal type_cast_4018_inst_ack_1 : boolean;
  signal if_stmt_4033_branch_req_0 : boolean;
  signal if_stmt_4033_branch_ack_1 : boolean;
  signal if_stmt_4033_branch_ack_0 : boolean;
  signal type_cast_4057_inst_req_0 : boolean;
  signal type_cast_4057_inst_ack_0 : boolean;
  signal type_cast_4057_inst_req_1 : boolean;
  signal type_cast_4057_inst_ack_1 : boolean;
  signal LOAD_col_high_4060_load_0_req_0 : boolean;
  signal LOAD_col_high_4060_load_0_ack_0 : boolean;
  signal LOAD_col_high_4060_load_0_req_1 : boolean;
  signal LOAD_col_high_4060_load_0_ack_1 : boolean;
  signal type_cast_4064_inst_req_0 : boolean;
  signal type_cast_4064_inst_ack_0 : boolean;
  signal type_cast_4064_inst_req_1 : boolean;
  signal type_cast_4064_inst_ack_1 : boolean;
  signal type_cast_4078_inst_req_0 : boolean;
  signal type_cast_4078_inst_ack_0 : boolean;
  signal type_cast_4078_inst_req_1 : boolean;
  signal type_cast_4078_inst_ack_1 : boolean;
  signal type_cast_4094_inst_req_0 : boolean;
  signal type_cast_4094_inst_ack_0 : boolean;
  signal type_cast_4094_inst_req_1 : boolean;
  signal type_cast_4094_inst_ack_1 : boolean;
  signal LOAD_row_high_4097_load_0_req_0 : boolean;
  signal LOAD_row_high_4097_load_0_ack_0 : boolean;
  signal LOAD_row_high_4097_load_0_req_1 : boolean;
  signal LOAD_row_high_4097_load_0_ack_1 : boolean;
  signal type_cast_4101_inst_req_0 : boolean;
  signal type_cast_4101_inst_ack_0 : boolean;
  signal type_cast_4101_inst_req_1 : boolean;
  signal type_cast_4101_inst_ack_1 : boolean;
  signal if_stmt_4125_branch_req_0 : boolean;
  signal if_stmt_4125_branch_ack_1 : boolean;
  signal if_stmt_4125_branch_ack_0 : boolean;
  signal LOAD_row_high_4156_load_0_req_0 : boolean;
  signal LOAD_row_high_4156_load_0_ack_0 : boolean;
  signal LOAD_row_high_4156_load_0_req_1 : boolean;
  signal LOAD_row_high_4156_load_0_ack_1 : boolean;
  signal type_cast_4160_inst_req_0 : boolean;
  signal type_cast_4160_inst_ack_0 : boolean;
  signal type_cast_4160_inst_req_1 : boolean;
  signal type_cast_4160_inst_ack_1 : boolean;
  signal LOAD_pad_4175_load_0_req_0 : boolean;
  signal LOAD_pad_4175_load_0_ack_0 : boolean;
  signal LOAD_pad_4175_load_0_req_1 : boolean;
  signal LOAD_pad_4175_load_0_ack_1 : boolean;
  signal LOAD_depth_high_4178_load_0_req_0 : boolean;
  signal LOAD_depth_high_4178_load_0_ack_0 : boolean;
  signal LOAD_depth_high_4178_load_0_req_1 : boolean;
  signal LOAD_depth_high_4178_load_0_ack_1 : boolean;
  signal ptr_deref_4550_load_0_ack_1 : boolean;
  signal ptr_deref_4550_load_0_req_1 : boolean;
  signal LOAD_col_high_4181_load_0_req_0 : boolean;
  signal type_cast_5037_inst_req_0 : boolean;
  signal LOAD_col_high_4181_load_0_ack_0 : boolean;
  signal type_cast_5037_inst_ack_0 : boolean;
  signal LOAD_col_high_4181_load_0_req_1 : boolean;
  signal LOAD_col_high_4181_load_0_ack_1 : boolean;
  signal array_obj_ref_5132_index_offset_ack_0 : boolean;
  signal if_stmt_4969_branch_ack_1 : boolean;
  signal type_cast_5037_inst_req_1 : boolean;
  signal type_cast_5037_inst_ack_1 : boolean;
  signal ptr_deref_4193_load_0_req_0 : boolean;
  signal ptr_deref_4193_load_0_ack_0 : boolean;
  signal ptr_deref_4193_load_0_req_1 : boolean;
  signal ptr_deref_4193_load_0_ack_1 : boolean;
  signal ptr_deref_5112_load_0_req_0 : boolean;
  signal ptr_deref_4205_load_0_req_0 : boolean;
  signal ptr_deref_4205_load_0_ack_0 : boolean;
  signal ptr_deref_5136_store_0_req_1 : boolean;
  signal ptr_deref_4205_load_0_req_1 : boolean;
  signal ptr_deref_4205_load_0_ack_1 : boolean;
  signal ptr_deref_5112_load_0_ack_0 : boolean;
  signal type_cast_4209_inst_req_0 : boolean;
  signal type_cast_4209_inst_ack_0 : boolean;
  signal type_cast_4209_inst_req_1 : boolean;
  signal type_cast_4209_inst_ack_1 : boolean;
  signal type_cast_4213_inst_req_0 : boolean;
  signal type_cast_4213_inst_ack_0 : boolean;
  signal if_stmt_4969_branch_ack_0 : boolean;
  signal type_cast_4213_inst_req_1 : boolean;
  signal type_cast_4213_inst_ack_1 : boolean;
  signal array_obj_ref_5024_index_offset_req_0 : boolean;
  signal type_cast_4252_inst_req_0 : boolean;
  signal type_cast_4252_inst_ack_0 : boolean;
  signal type_cast_4252_inst_req_1 : boolean;
  signal type_cast_4252_inst_ack_1 : boolean;
  signal array_obj_ref_5024_index_offset_ack_0 : boolean;
  signal type_cast_4321_inst_req_0 : boolean;
  signal type_cast_4321_inst_ack_0 : boolean;
  signal type_cast_4321_inst_req_1 : boolean;
  signal type_cast_4321_inst_ack_1 : boolean;
  signal if_stmt_4330_branch_req_0 : boolean;
  signal if_stmt_4330_branch_ack_1 : boolean;
  signal if_stmt_4330_branch_ack_0 : boolean;
  signal ptr_deref_5112_load_0_req_1 : boolean;
  signal array_obj_ref_5132_index_offset_req_1 : boolean;
  signal LOAD_row_high_4338_load_0_req_0 : boolean;
  signal type_cast_5101_inst_req_0 : boolean;
  signal LOAD_row_high_4338_load_0_ack_0 : boolean;
  signal type_cast_5101_inst_ack_0 : boolean;
  signal ptr_deref_5136_store_0_ack_1 : boolean;
  signal LOAD_row_high_4338_load_0_req_1 : boolean;
  signal LOAD_row_high_4338_load_0_ack_1 : boolean;
  signal ptr_deref_5112_load_0_ack_1 : boolean;
  signal type_cast_5101_inst_req_1 : boolean;
  signal array_obj_ref_5024_index_offset_req_1 : boolean;
  signal array_obj_ref_5132_index_offset_ack_1 : boolean;
  signal type_cast_4342_inst_req_0 : boolean;
  signal type_cast_4342_inst_ack_0 : boolean;
  signal type_cast_4342_inst_req_1 : boolean;
  signal type_cast_5101_inst_ack_1 : boolean;
  signal type_cast_4342_inst_ack_1 : boolean;
  signal array_obj_ref_5024_index_offset_ack_1 : boolean;
  signal if_stmt_4356_branch_req_0 : boolean;
  signal if_stmt_4356_branch_ack_1 : boolean;
  signal if_stmt_4356_branch_ack_0 : boolean;
  signal addr_of_5108_final_reg_req_0 : boolean;
  signal type_cast_4366_inst_req_0 : boolean;
  signal type_cast_4366_inst_ack_0 : boolean;
  signal type_cast_4366_inst_req_1 : boolean;
  signal type_cast_4366_inst_ack_1 : boolean;
  signal addr_of_5108_final_reg_ack_0 : boolean;
  signal if_stmt_4375_branch_req_0 : boolean;
  signal if_stmt_4375_branch_ack_1 : boolean;
  signal if_stmt_4375_branch_ack_0 : boolean;
  signal LOAD_col_high_4383_load_0_req_0 : boolean;
  signal LOAD_col_high_4383_load_0_ack_0 : boolean;
  signal LOAD_col_high_4383_load_0_req_1 : boolean;
  signal LOAD_col_high_4383_load_0_ack_1 : boolean;
  signal type_cast_4387_inst_req_0 : boolean;
  signal type_cast_4387_inst_ack_0 : boolean;
  signal type_cast_4387_inst_req_1 : boolean;
  signal type_cast_4387_inst_ack_1 : boolean;
  signal if_stmt_4407_branch_req_0 : boolean;
  signal if_stmt_4407_branch_ack_1 : boolean;
  signal if_stmt_4407_branch_ack_0 : boolean;
  signal type_cast_4417_inst_req_0 : boolean;
  signal type_cast_4417_inst_ack_0 : boolean;
  signal type_cast_4417_inst_req_1 : boolean;
  signal type_cast_4417_inst_ack_1 : boolean;
  signal type_cast_4422_inst_req_0 : boolean;
  signal type_cast_4422_inst_ack_0 : boolean;
  signal type_cast_4422_inst_req_1 : boolean;
  signal type_cast_4422_inst_ack_1 : boolean;
  signal type_cast_4456_inst_req_0 : boolean;
  signal type_cast_4456_inst_ack_0 : boolean;
  signal type_cast_4456_inst_req_1 : boolean;
  signal type_cast_4456_inst_ack_1 : boolean;
  signal array_obj_ref_4462_index_offset_req_0 : boolean;
  signal array_obj_ref_4462_index_offset_ack_0 : boolean;
  signal array_obj_ref_4462_index_offset_req_1 : boolean;
  signal array_obj_ref_4462_index_offset_ack_1 : boolean;
  signal addr_of_4463_final_reg_req_0 : boolean;
  signal addr_of_4463_final_reg_ack_0 : boolean;
  signal addr_of_4463_final_reg_req_1 : boolean;
  signal addr_of_4463_final_reg_ack_1 : boolean;
  signal ptr_deref_4466_store_0_req_0 : boolean;
  signal ptr_deref_4466_store_0_ack_0 : boolean;
  signal ptr_deref_4466_store_0_req_1 : boolean;
  signal ptr_deref_4466_store_0_ack_1 : boolean;
  signal type_cast_4475_inst_req_0 : boolean;
  signal type_cast_4475_inst_ack_0 : boolean;
  signal type_cast_4475_inst_req_1 : boolean;
  signal type_cast_4475_inst_ack_1 : boolean;
  signal type_cast_4539_inst_req_0 : boolean;
  signal type_cast_4539_inst_ack_0 : boolean;
  signal type_cast_4539_inst_req_1 : boolean;
  signal type_cast_4539_inst_ack_1 : boolean;
  signal array_obj_ref_4545_index_offset_req_0 : boolean;
  signal array_obj_ref_4545_index_offset_ack_0 : boolean;
  signal array_obj_ref_4545_index_offset_req_1 : boolean;
  signal array_obj_ref_4545_index_offset_ack_1 : boolean;
  signal addr_of_4546_final_reg_req_0 : boolean;
  signal addr_of_4546_final_reg_ack_0 : boolean;
  signal addr_of_4546_final_reg_req_1 : boolean;
  signal addr_of_4546_final_reg_ack_1 : boolean;
  signal type_cast_4582_inst_req_1 : boolean;
  signal type_cast_4582_inst_ack_1 : boolean;
  signal if_stmt_4597_branch_req_0 : boolean;
  signal if_stmt_4597_branch_ack_1 : boolean;
  signal if_stmt_4597_branch_ack_0 : boolean;
  signal type_cast_4621_inst_req_0 : boolean;
  signal type_cast_4621_inst_ack_0 : boolean;
  signal type_cast_4621_inst_req_1 : boolean;
  signal type_cast_4621_inst_ack_1 : boolean;
  signal LOAD_col_high_4624_load_0_req_0 : boolean;
  signal LOAD_col_high_4624_load_0_ack_0 : boolean;
  signal LOAD_col_high_4624_load_0_req_1 : boolean;
  signal LOAD_col_high_4624_load_0_ack_1 : boolean;
  signal type_cast_4628_inst_req_0 : boolean;
  signal type_cast_4628_inst_ack_0 : boolean;
  signal type_cast_4628_inst_req_1 : boolean;
  signal type_cast_4628_inst_ack_1 : boolean;
  signal type_cast_4648_inst_req_0 : boolean;
  signal type_cast_4648_inst_ack_0 : boolean;
  signal type_cast_4648_inst_req_1 : boolean;
  signal type_cast_4648_inst_ack_1 : boolean;
  signal type_cast_4665_inst_req_0 : boolean;
  signal type_cast_4665_inst_ack_0 : boolean;
  signal type_cast_4665_inst_req_1 : boolean;
  signal type_cast_4665_inst_ack_1 : boolean;
  signal LOAD_row_high_4668_load_0_req_0 : boolean;
  signal LOAD_row_high_4668_load_0_ack_0 : boolean;
  signal LOAD_row_high_4668_load_0_req_1 : boolean;
  signal LOAD_row_high_4668_load_0_ack_1 : boolean;
  signal type_cast_4672_inst_req_0 : boolean;
  signal type_cast_4672_inst_ack_0 : boolean;
  signal type_cast_4672_inst_req_1 : boolean;
  signal type_cast_4672_inst_ack_1 : boolean;
  signal if_stmt_4684_branch_req_0 : boolean;
  signal if_stmt_4684_branch_ack_1 : boolean;
  signal if_stmt_4684_branch_ack_0 : boolean;
  signal LOAD_col_high_4715_load_0_req_0 : boolean;
  signal LOAD_col_high_4715_load_0_ack_0 : boolean;
  signal LOAD_col_high_4715_load_0_req_1 : boolean;
  signal LOAD_col_high_4715_load_0_ack_1 : boolean;
  signal type_cast_4719_inst_req_0 : boolean;
  signal type_cast_4719_inst_ack_0 : boolean;
  signal type_cast_4719_inst_req_1 : boolean;
  signal type_cast_4719_inst_ack_1 : boolean;
  signal LOAD_row_high_4728_load_0_req_0 : boolean;
  signal LOAD_row_high_4728_load_0_ack_0 : boolean;
  signal LOAD_row_high_4728_load_0_req_1 : boolean;
  signal LOAD_row_high_4728_load_0_ack_1 : boolean;
  signal type_cast_4732_inst_req_0 : boolean;
  signal type_cast_4732_inst_ack_0 : boolean;
  signal type_cast_4732_inst_req_1 : boolean;
  signal type_cast_4732_inst_ack_1 : boolean;
  signal LOAD_pad_4747_load_0_req_0 : boolean;
  signal LOAD_pad_4747_load_0_ack_0 : boolean;
  signal LOAD_pad_4747_load_0_req_1 : boolean;
  signal LOAD_pad_4747_load_0_ack_1 : boolean;
  signal type_cast_5018_inst_ack_1 : boolean;
  signal type_cast_5018_inst_req_1 : boolean;
  signal LOAD_depth_high_4750_load_0_req_0 : boolean;
  signal LOAD_depth_high_4750_load_0_ack_0 : boolean;
  signal type_cast_5018_inst_ack_0 : boolean;
  signal LOAD_depth_high_4750_load_0_req_1 : boolean;
  signal LOAD_depth_high_4750_load_0_ack_1 : boolean;
  signal type_cast_5018_inst_req_0 : boolean;
  signal ptr_deref_4762_load_0_req_0 : boolean;
  signal ptr_deref_4762_load_0_ack_0 : boolean;
  signal ptr_deref_4762_load_0_req_1 : boolean;
  signal ptr_deref_4762_load_0_ack_1 : boolean;
  signal array_obj_ref_5132_index_offset_req_0 : boolean;
  signal type_cast_5126_inst_ack_1 : boolean;
  signal type_cast_5126_inst_req_1 : boolean;
  signal type_cast_5126_inst_ack_0 : boolean;
  signal type_cast_4984_inst_ack_1 : boolean;
  signal type_cast_4984_inst_req_1 : boolean;
  signal addr_of_5025_final_reg_ack_1 : boolean;
  signal addr_of_5025_final_reg_req_1 : boolean;
  signal ptr_deref_4774_load_0_req_0 : boolean;
  signal ptr_deref_5028_store_0_ack_1 : boolean;
  signal ptr_deref_4774_load_0_ack_0 : boolean;
  signal ptr_deref_4774_load_0_req_1 : boolean;
  signal ptr_deref_5028_store_0_req_1 : boolean;
  signal ptr_deref_4774_load_0_ack_1 : boolean;
  signal type_cast_4984_inst_ack_0 : boolean;
  signal type_cast_4984_inst_req_0 : boolean;
  signal type_cast_5126_inst_req_0 : boolean;
  signal type_cast_4778_inst_req_0 : boolean;
  signal type_cast_4778_inst_ack_0 : boolean;
  signal array_obj_ref_5107_index_offset_ack_1 : boolean;
  signal type_cast_4778_inst_req_1 : boolean;
  signal type_cast_4778_inst_ack_1 : boolean;
  signal type_cast_5144_inst_ack_1 : boolean;
  signal type_cast_5144_inst_req_1 : boolean;
  signal if_stmt_4969_branch_req_0 : boolean;
  signal type_cast_4782_inst_req_0 : boolean;
  signal type_cast_4782_inst_ack_0 : boolean;
  signal array_obj_ref_5107_index_offset_req_1 : boolean;
  signal type_cast_4782_inst_req_1 : boolean;
  signal type_cast_4782_inst_ack_1 : boolean;
  signal type_cast_4821_inst_req_0 : boolean;
  signal type_cast_4821_inst_ack_0 : boolean;
  signal type_cast_4821_inst_req_1 : boolean;
  signal type_cast_4821_inst_ack_1 : boolean;
  signal type_cast_5144_inst_ack_0 : boolean;
  signal type_cast_5144_inst_req_0 : boolean;
  signal type_cast_4889_inst_req_0 : boolean;
  signal type_cast_4889_inst_ack_0 : boolean;
  signal type_cast_4889_inst_req_1 : boolean;
  signal type_cast_4889_inst_ack_1 : boolean;
  signal array_obj_ref_5107_index_offset_ack_0 : boolean;
  signal if_stmt_4898_branch_req_0 : boolean;
  signal ptr_deref_5028_store_0_ack_0 : boolean;
  signal array_obj_ref_5107_index_offset_req_0 : boolean;
  signal if_stmt_4898_branch_ack_1 : boolean;
  signal if_stmt_4898_branch_ack_0 : boolean;
  signal ptr_deref_5028_store_0_req_0 : boolean;
  signal addr_of_5025_final_reg_ack_0 : boolean;
  signal LOAD_row_high_4906_load_0_req_0 : boolean;
  signal LOAD_row_high_4906_load_0_ack_0 : boolean;
  signal addr_of_5025_final_reg_req_0 : boolean;
  signal LOAD_row_high_4906_load_0_req_1 : boolean;
  signal LOAD_row_high_4906_load_0_ack_1 : boolean;
  signal ptr_deref_5136_store_0_ack_0 : boolean;
  signal ptr_deref_5136_store_0_req_0 : boolean;
  signal addr_of_5133_final_reg_ack_1 : boolean;
  signal addr_of_5133_final_reg_req_1 : boolean;
  signal type_cast_4910_inst_req_0 : boolean;
  signal type_cast_4910_inst_ack_0 : boolean;
  signal type_cast_4910_inst_req_1 : boolean;
  signal addr_of_5108_final_reg_ack_1 : boolean;
  signal type_cast_4910_inst_ack_1 : boolean;
  signal type_cast_4979_inst_ack_1 : boolean;
  signal addr_of_5133_final_reg_ack_0 : boolean;
  signal if_stmt_4924_branch_req_0 : boolean;
  signal type_cast_4979_inst_req_1 : boolean;
  signal if_stmt_4924_branch_ack_1 : boolean;
  signal if_stmt_4924_branch_ack_0 : boolean;
  signal addr_of_5133_final_reg_req_0 : boolean;
  signal type_cast_4934_inst_req_0 : boolean;
  signal addr_of_5108_final_reg_req_1 : boolean;
  signal type_cast_4934_inst_ack_0 : boolean;
  signal type_cast_4934_inst_req_1 : boolean;
  signal type_cast_4934_inst_ack_1 : boolean;
  signal type_cast_4979_inst_ack_0 : boolean;
  signal if_stmt_4943_branch_req_0 : boolean;
  signal type_cast_4979_inst_req_0 : boolean;
  signal if_stmt_4943_branch_ack_1 : boolean;
  signal if_stmt_4943_branch_ack_0 : boolean;
  signal LOAD_col_high_4951_load_0_req_0 : boolean;
  signal LOAD_col_high_4951_load_0_ack_0 : boolean;
  signal LOAD_col_high_4951_load_0_req_1 : boolean;
  signal LOAD_col_high_4951_load_0_ack_1 : boolean;
  signal type_cast_2437_inst_ack_1 : boolean;
  signal type_cast_2602_inst_req_0 : boolean;
  signal type_cast_4955_inst_req_0 : boolean;
  signal type_cast_4955_inst_ack_0 : boolean;
  signal type_cast_4955_inst_req_1 : boolean;
  signal type_cast_4955_inst_ack_1 : boolean;
  signal if_stmt_5159_branch_req_0 : boolean;
  signal if_stmt_5159_branch_ack_1 : boolean;
  signal if_stmt_5159_branch_ack_0 : boolean;
  signal type_cast_5183_inst_req_0 : boolean;
  signal type_cast_5183_inst_ack_0 : boolean;
  signal type_cast_5183_inst_req_1 : boolean;
  signal type_cast_5183_inst_ack_1 : boolean;
  signal LOAD_col_high_5186_load_0_req_0 : boolean;
  signal LOAD_col_high_5186_load_0_ack_0 : boolean;
  signal LOAD_col_high_5186_load_0_req_1 : boolean;
  signal LOAD_col_high_5186_load_0_ack_1 : boolean;
  signal type_cast_5190_inst_req_0 : boolean;
  signal type_cast_5190_inst_ack_0 : boolean;
  signal type_cast_5190_inst_req_1 : boolean;
  signal type_cast_5190_inst_ack_1 : boolean;
  signal type_cast_5204_inst_req_0 : boolean;
  signal type_cast_5204_inst_ack_0 : boolean;
  signal type_cast_5204_inst_req_1 : boolean;
  signal type_cast_5204_inst_ack_1 : boolean;
  signal type_cast_5220_inst_req_0 : boolean;
  signal type_cast_5220_inst_ack_0 : boolean;
  signal type_cast_5220_inst_req_1 : boolean;
  signal type_cast_5220_inst_ack_1 : boolean;
  signal LOAD_row_high_5223_load_0_req_0 : boolean;
  signal LOAD_row_high_5223_load_0_ack_0 : boolean;
  signal LOAD_row_high_5223_load_0_req_1 : boolean;
  signal LOAD_row_high_5223_load_0_ack_1 : boolean;
  signal type_cast_2437_inst_req_1 : boolean;
  signal type_cast_2596_inst_req_0 : boolean;
  signal type_cast_2437_inst_ack_0 : boolean;
  signal type_cast_5227_inst_req_0 : boolean;
  signal type_cast_2437_inst_req_0 : boolean;
  signal type_cast_5227_inst_ack_0 : boolean;
  signal type_cast_5227_inst_req_1 : boolean;
  signal type_cast_5227_inst_ack_1 : boolean;
  signal if_stmt_5239_branch_req_0 : boolean;
  signal if_stmt_5239_branch_ack_1 : boolean;
  signal phi_stmt_2421_req_0 : boolean;
  signal if_stmt_5239_branch_ack_0 : boolean;
  signal type_cast_2424_inst_ack_1 : boolean;
  signal type_cast_2424_inst_req_1 : boolean;
  signal call_stmt_5270_call_req_0 : boolean;
  signal call_stmt_5270_call_ack_0 : boolean;
  signal call_stmt_5270_call_req_1 : boolean;
  signal call_stmt_5270_call_ack_1 : boolean;
  signal phi_stmt_2597_req_1 : boolean;
  signal phi_stmt_2434_req_0 : boolean;
  signal phi_stmt_899_req_0 : boolean;
  signal phi_stmt_906_req_0 : boolean;
  signal phi_stmt_913_req_0 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal phi_stmt_899_req_1 : boolean;
  signal type_cast_912_inst_req_0 : boolean;
  signal type_cast_912_inst_ack_0 : boolean;
  signal type_cast_912_inst_req_1 : boolean;
  signal type_cast_912_inst_ack_1 : boolean;
  signal phi_stmt_906_req_1 : boolean;
  signal phi_stmt_2428_req_0 : boolean;
  signal type_cast_2433_inst_ack_0 : boolean;
  signal type_cast_919_inst_req_0 : boolean;
  signal type_cast_2431_inst_ack_1 : boolean;
  signal type_cast_919_inst_ack_0 : boolean;
  signal type_cast_919_inst_req_1 : boolean;
  signal phi_stmt_2434_req_1 : boolean;
  signal type_cast_919_inst_ack_1 : boolean;
  signal phi_stmt_913_req_1 : boolean;
  signal type_cast_2439_inst_ack_1 : boolean;
  signal type_cast_2431_inst_req_1 : boolean;
  signal type_cast_2602_inst_ack_1 : boolean;
  signal phi_stmt_899_ack_0 : boolean;
  signal phi_stmt_906_ack_0 : boolean;
  signal phi_stmt_913_ack_0 : boolean;
  signal type_cast_2433_inst_req_0 : boolean;
  signal type_cast_2439_inst_req_1 : boolean;
  signal phi_stmt_2434_ack_0 : boolean;
  signal phi_stmt_2421_req_1 : boolean;
  signal type_cast_2424_inst_ack_0 : boolean;
  signal type_cast_2424_inst_req_0 : boolean;
  signal type_cast_2431_inst_ack_0 : boolean;
  signal type_cast_2431_inst_req_0 : boolean;
  signal type_cast_2439_inst_ack_0 : boolean;
  signal type_cast_2602_inst_req_1 : boolean;
  signal type_cast_2439_inst_req_0 : boolean;
  signal phi_stmt_2428_ack_0 : boolean;
  signal type_cast_2602_inst_ack_0 : boolean;
  signal phi_stmt_2421_ack_0 : boolean;
  signal type_cast_1318_inst_req_0 : boolean;
  signal type_cast_1318_inst_ack_0 : boolean;
  signal type_cast_1318_inst_req_1 : boolean;
  signal phi_stmt_2428_req_1 : boolean;
  signal type_cast_1318_inst_ack_1 : boolean;
  signal phi_stmt_1313_req_1 : boolean;
  signal phi_stmt_1319_req_0 : boolean;
  signal phi_stmt_2590_req_1 : boolean;
  signal type_cast_2596_inst_ack_1 : boolean;
  signal type_cast_2596_inst_req_1 : boolean;
  signal type_cast_1310_inst_req_0 : boolean;
  signal type_cast_1310_inst_ack_0 : boolean;
  signal type_cast_2433_inst_ack_1 : boolean;
  signal type_cast_1310_inst_req_1 : boolean;
  signal type_cast_2433_inst_req_1 : boolean;
  signal type_cast_1310_inst_ack_1 : boolean;
  signal phi_stmt_1307_req_0 : boolean;
  signal type_cast_2596_inst_ack_0 : boolean;
  signal type_cast_1316_inst_req_0 : boolean;
  signal type_cast_1316_inst_ack_0 : boolean;
  signal type_cast_1316_inst_req_1 : boolean;
  signal type_cast_1316_inst_ack_1 : boolean;
  signal phi_stmt_1313_req_0 : boolean;
  signal type_cast_1325_inst_req_0 : boolean;
  signal type_cast_1325_inst_ack_0 : boolean;
  signal type_cast_1325_inst_req_1 : boolean;
  signal type_cast_1325_inst_ack_1 : boolean;
  signal phi_stmt_1319_req_1 : boolean;
  signal type_cast_1312_inst_req_0 : boolean;
  signal type_cast_1312_inst_ack_0 : boolean;
  signal type_cast_1312_inst_req_1 : boolean;
  signal type_cast_1312_inst_ack_1 : boolean;
  signal phi_stmt_1307_req_1 : boolean;
  signal phi_stmt_1307_ack_0 : boolean;
  signal phi_stmt_1313_ack_0 : boolean;
  signal phi_stmt_1319_ack_0 : boolean;
  signal type_cast_4142_inst_req_1 : boolean;
  signal type_cast_1468_inst_req_0 : boolean;
  signal type_cast_1468_inst_ack_0 : boolean;
  signal type_cast_4303_inst_req_0 : boolean;
  signal type_cast_1468_inst_req_1 : boolean;
  signal type_cast_1468_inst_ack_1 : boolean;
  signal phi_stmt_1463_req_1 : boolean;
  signal type_cast_4142_inst_ack_1 : boolean;
  signal type_cast_1475_inst_req_0 : boolean;
  signal type_cast_1475_inst_ack_0 : boolean;
  signal type_cast_1475_inst_req_1 : boolean;
  signal type_cast_1475_inst_ack_1 : boolean;
  signal phi_stmt_1469_req_1 : boolean;
  signal type_cast_1482_inst_req_0 : boolean;
  signal type_cast_1482_inst_ack_0 : boolean;
  signal type_cast_1482_inst_req_1 : boolean;
  signal type_cast_1482_inst_ack_1 : boolean;
  signal phi_stmt_1476_req_1 : boolean;
  signal type_cast_4303_inst_ack_0 : boolean;
  signal type_cast_1466_inst_req_0 : boolean;
  signal type_cast_1466_inst_ack_0 : boolean;
  signal type_cast_1466_inst_req_1 : boolean;
  signal type_cast_1466_inst_ack_1 : boolean;
  signal phi_stmt_1463_req_0 : boolean;
  signal phi_stmt_1469_req_0 : boolean;
  signal phi_stmt_1476_req_0 : boolean;
  signal phi_stmt_4139_req_0 : boolean;
  signal type_cast_4303_inst_req_1 : boolean;
  signal type_cast_4303_inst_ack_1 : boolean;
  signal phi_stmt_1463_ack_0 : boolean;
  signal phi_stmt_1469_ack_0 : boolean;
  signal phi_stmt_1476_ack_0 : boolean;
  signal phi_stmt_4297_req_1 : boolean;
  signal type_cast_4316_inst_req_0 : boolean;
  signal type_cast_4316_inst_ack_0 : boolean;
  signal phi_stmt_1868_req_1 : boolean;
  signal type_cast_1867_inst_req_0 : boolean;
  signal type_cast_1867_inst_ack_0 : boolean;
  signal type_cast_1867_inst_req_1 : boolean;
  signal type_cast_1867_inst_ack_1 : boolean;
  signal phi_stmt_1862_req_1 : boolean;
  signal type_cast_1861_inst_req_0 : boolean;
  signal type_cast_1861_inst_ack_0 : boolean;
  signal type_cast_1861_inst_req_1 : boolean;
  signal type_cast_1861_inst_ack_1 : boolean;
  signal phi_stmt_1856_req_1 : boolean;
  signal type_cast_1871_inst_req_0 : boolean;
  signal type_cast_1871_inst_ack_0 : boolean;
  signal type_cast_1871_inst_req_1 : boolean;
  signal type_cast_1871_inst_ack_1 : boolean;
  signal phi_stmt_1868_req_0 : boolean;
  signal type_cast_1865_inst_req_0 : boolean;
  signal type_cast_1865_inst_ack_0 : boolean;
  signal type_cast_1865_inst_req_1 : boolean;
  signal type_cast_1865_inst_ack_1 : boolean;
  signal phi_stmt_1862_req_0 : boolean;
  signal type_cast_1859_inst_req_0 : boolean;
  signal type_cast_1859_inst_ack_0 : boolean;
  signal type_cast_1859_inst_req_1 : boolean;
  signal type_cast_1859_inst_ack_1 : boolean;
  signal phi_stmt_1856_req_0 : boolean;
  signal phi_stmt_1856_ack_0 : boolean;
  signal phi_stmt_1862_ack_0 : boolean;
  signal phi_stmt_1868_ack_0 : boolean;
  signal type_cast_2018_inst_req_0 : boolean;
  signal type_cast_2018_inst_ack_0 : boolean;
  signal type_cast_2018_inst_req_1 : boolean;
  signal type_cast_2018_inst_ack_1 : boolean;
  signal phi_stmt_2015_req_0 : boolean;
  signal type_cast_2031_inst_req_0 : boolean;
  signal type_cast_2031_inst_ack_0 : boolean;
  signal type_cast_2031_inst_req_1 : boolean;
  signal type_cast_2031_inst_ack_1 : boolean;
  signal phi_stmt_2028_req_0 : boolean;
  signal type_cast_2027_inst_req_0 : boolean;
  signal type_cast_2027_inst_ack_0 : boolean;
  signal type_cast_2027_inst_req_1 : boolean;
  signal type_cast_2027_inst_ack_1 : boolean;
  signal phi_stmt_2022_req_1 : boolean;
  signal phi_stmt_2015_req_1 : boolean;
  signal phi_stmt_2028_req_1 : boolean;
  signal type_cast_2025_inst_req_0 : boolean;
  signal type_cast_2025_inst_ack_0 : boolean;
  signal type_cast_2025_inst_req_1 : boolean;
  signal type_cast_2025_inst_ack_1 : boolean;
  signal phi_stmt_2022_req_0 : boolean;
  signal phi_stmt_2015_ack_0 : boolean;
  signal phi_stmt_2022_ack_0 : boolean;
  signal phi_stmt_2028_ack_0 : boolean;
  signal type_cast_2608_inst_req_0 : boolean;
  signal type_cast_2608_inst_ack_0 : boolean;
  signal type_cast_2608_inst_req_1 : boolean;
  signal type_cast_2608_inst_ack_1 : boolean;
  signal phi_stmt_2603_req_1 : boolean;
  signal phi_stmt_2590_req_0 : boolean;
  signal type_cast_2600_inst_req_0 : boolean;
  signal type_cast_2600_inst_ack_0 : boolean;
  signal type_cast_2600_inst_req_1 : boolean;
  signal type_cast_2600_inst_ack_1 : boolean;
  signal phi_stmt_2597_req_0 : boolean;
  signal type_cast_2606_inst_req_0 : boolean;
  signal type_cast_2606_inst_ack_0 : boolean;
  signal type_cast_2606_inst_req_1 : boolean;
  signal type_cast_2606_inst_ack_1 : boolean;
  signal phi_stmt_2603_req_0 : boolean;
  signal phi_stmt_2590_ack_0 : boolean;
  signal phi_stmt_2597_ack_0 : boolean;
  signal phi_stmt_2603_ack_0 : boolean;
  signal phi_stmt_2982_req_1 : boolean;
  signal type_cast_2994_inst_req_0 : boolean;
  signal type_cast_2994_inst_ack_0 : boolean;
  signal type_cast_2994_inst_req_1 : boolean;
  signal type_cast_2994_inst_ack_1 : boolean;
  signal phi_stmt_2989_req_1 : boolean;
  signal type_cast_3000_inst_req_0 : boolean;
  signal type_cast_3000_inst_ack_0 : boolean;
  signal type_cast_3000_inst_req_1 : boolean;
  signal type_cast_3000_inst_ack_1 : boolean;
  signal phi_stmt_2995_req_1 : boolean;
  signal type_cast_2985_inst_req_0 : boolean;
  signal type_cast_2985_inst_ack_0 : boolean;
  signal type_cast_2985_inst_req_1 : boolean;
  signal type_cast_2985_inst_ack_1 : boolean;
  signal phi_stmt_2982_req_0 : boolean;
  signal type_cast_2992_inst_req_0 : boolean;
  signal type_cast_2992_inst_ack_0 : boolean;
  signal type_cast_2992_inst_req_1 : boolean;
  signal type_cast_2992_inst_ack_1 : boolean;
  signal phi_stmt_2989_req_0 : boolean;
  signal type_cast_2998_inst_req_0 : boolean;
  signal type_cast_2998_inst_ack_0 : boolean;
  signal type_cast_2998_inst_req_1 : boolean;
  signal type_cast_2998_inst_ack_1 : boolean;
  signal phi_stmt_2995_req_0 : boolean;
  signal phi_stmt_2982_ack_0 : boolean;
  signal phi_stmt_2989_ack_0 : boolean;
  signal phi_stmt_2995_ack_0 : boolean;
  signal type_cast_3157_inst_req_0 : boolean;
  signal type_cast_3157_inst_ack_0 : boolean;
  signal type_cast_3157_inst_req_1 : boolean;
  signal type_cast_3157_inst_ack_1 : boolean;
  signal phi_stmt_3154_req_0 : boolean;
  signal type_cast_3153_inst_req_0 : boolean;
  signal type_cast_3153_inst_ack_0 : boolean;
  signal type_cast_3153_inst_req_1 : boolean;
  signal type_cast_3153_inst_ack_1 : boolean;
  signal phi_stmt_3148_req_1 : boolean;
  signal type_cast_3144_inst_req_0 : boolean;
  signal type_cast_3144_inst_ack_0 : boolean;
  signal type_cast_3144_inst_req_1 : boolean;
  signal type_cast_3144_inst_ack_1 : boolean;
  signal phi_stmt_3141_req_0 : boolean;
  signal phi_stmt_3154_req_1 : boolean;
  signal type_cast_3151_inst_req_0 : boolean;
  signal type_cast_3151_inst_ack_0 : boolean;
  signal type_cast_3151_inst_req_1 : boolean;
  signal type_cast_3151_inst_ack_1 : boolean;
  signal phi_stmt_3148_req_0 : boolean;
  signal phi_stmt_3141_req_1 : boolean;
  signal phi_stmt_3141_ack_0 : boolean;
  signal phi_stmt_3148_ack_0 : boolean;
  signal phi_stmt_3154_ack_0 : boolean;
  signal phi_stmt_4139_ack_0 : boolean;
  signal phi_stmt_4132_ack_0 : boolean;
  signal type_cast_4709_inst_ack_1 : boolean;
  signal phi_stmt_4698_req_1 : boolean;
  signal phi_stmt_4145_req_0 : boolean;
  signal type_cast_4148_inst_ack_1 : boolean;
  signal type_cast_4148_inst_req_1 : boolean;
  signal phi_stmt_3559_req_1 : boolean;
  signal type_cast_4148_inst_ack_0 : boolean;
  signal type_cast_4148_inst_req_0 : boolean;
  signal type_cast_3571_inst_req_0 : boolean;
  signal type_cast_3571_inst_ack_0 : boolean;
  signal type_cast_3571_inst_req_1 : boolean;
  signal phi_stmt_4310_ack_0 : boolean;
  signal type_cast_3571_inst_ack_1 : boolean;
  signal phi_stmt_3566_req_1 : boolean;
  signal type_cast_3575_inst_req_0 : boolean;
  signal type_cast_3575_inst_ack_0 : boolean;
  signal phi_stmt_4304_ack_0 : boolean;
  signal type_cast_3575_inst_req_1 : boolean;
  signal phi_stmt_4297_ack_0 : boolean;
  signal type_cast_3575_inst_ack_1 : boolean;
  signal phi_stmt_3572_req_0 : boolean;
  signal type_cast_4709_inst_req_1 : boolean;
  signal phi_stmt_4704_req_0 : boolean;
  signal type_cast_4707_inst_ack_1 : boolean;
  signal type_cast_3562_inst_req_0 : boolean;
  signal type_cast_3562_inst_ack_0 : boolean;
  signal type_cast_3562_inst_req_1 : boolean;
  signal phi_stmt_4310_req_0 : boolean;
  signal type_cast_3562_inst_ack_1 : boolean;
  signal phi_stmt_3559_req_0 : boolean;
  signal type_cast_4707_inst_req_1 : boolean;
  signal type_cast_3569_inst_req_0 : boolean;
  signal type_cast_3569_inst_ack_0 : boolean;
  signal type_cast_3569_inst_req_1 : boolean;
  signal type_cast_3569_inst_ack_1 : boolean;
  signal phi_stmt_3566_req_0 : boolean;
  signal type_cast_4142_inst_ack_0 : boolean;
  signal type_cast_4707_inst_ack_0 : boolean;
  signal type_cast_3577_inst_req_0 : boolean;
  signal type_cast_3577_inst_ack_0 : boolean;
  signal type_cast_3577_inst_req_1 : boolean;
  signal type_cast_3577_inst_ack_1 : boolean;
  signal phi_stmt_3572_req_1 : boolean;
  signal type_cast_4707_inst_req_0 : boolean;
  signal type_cast_4701_inst_ack_0 : boolean;
  signal phi_stmt_3559_ack_0 : boolean;
  signal phi_stmt_3566_ack_0 : boolean;
  signal phi_stmt_3572_ack_0 : boolean;
  signal phi_stmt_4304_req_0 : boolean;
  signal type_cast_4307_inst_ack_1 : boolean;
  signal type_cast_4703_inst_ack_1 : boolean;
  signal phi_stmt_4304_req_1 : boolean;
  signal type_cast_3731_inst_req_0 : boolean;
  signal type_cast_3731_inst_ack_0 : boolean;
  signal type_cast_4307_inst_req_1 : boolean;
  signal type_cast_3731_inst_req_1 : boolean;
  signal type_cast_3731_inst_ack_1 : boolean;
  signal phi_stmt_3728_req_0 : boolean;
  signal type_cast_3740_inst_req_0 : boolean;
  signal type_cast_3740_inst_ack_0 : boolean;
  signal type_cast_3740_inst_req_1 : boolean;
  signal type_cast_3740_inst_ack_1 : boolean;
  signal phi_stmt_3735_req_1 : boolean;
  signal type_cast_4309_inst_ack_1 : boolean;
  signal type_cast_3744_inst_req_0 : boolean;
  signal type_cast_3744_inst_ack_0 : boolean;
  signal type_cast_3744_inst_req_1 : boolean;
  signal type_cast_3744_inst_ack_1 : boolean;
  signal phi_stmt_3741_req_0 : boolean;
  signal type_cast_4307_inst_ack_0 : boolean;
  signal type_cast_4709_inst_ack_0 : boolean;
  signal phi_stmt_3728_req_1 : boolean;
  signal type_cast_4309_inst_req_1 : boolean;
  signal type_cast_3738_inst_req_0 : boolean;
  signal type_cast_3738_inst_ack_0 : boolean;
  signal type_cast_4307_inst_req_0 : boolean;
  signal type_cast_3738_inst_req_1 : boolean;
  signal type_cast_3738_inst_ack_1 : boolean;
  signal phi_stmt_3735_req_0 : boolean;
  signal type_cast_4142_inst_req_0 : boolean;
  signal type_cast_3746_inst_req_0 : boolean;
  signal type_cast_3746_inst_ack_0 : boolean;
  signal type_cast_3746_inst_req_1 : boolean;
  signal type_cast_3746_inst_ack_1 : boolean;
  signal phi_stmt_3741_req_1 : boolean;
  signal type_cast_4701_inst_req_0 : boolean;
  signal phi_stmt_3728_ack_0 : boolean;
  signal phi_stmt_3735_ack_0 : boolean;
  signal phi_stmt_3741_ack_0 : boolean;
  signal type_cast_4703_inst_req_1 : boolean;
  signal type_cast_4703_inst_ack_0 : boolean;
  signal phi_stmt_4297_req_0 : boolean;
  signal type_cast_4703_inst_req_0 : boolean;
  signal phi_stmt_4691_req_1 : boolean;
  signal type_cast_4309_inst_ack_0 : boolean;
  signal type_cast_4709_inst_req_0 : boolean;
  signal type_cast_4309_inst_req_0 : boolean;
  signal phi_stmt_4310_req_1 : boolean;
  signal type_cast_4316_inst_ack_1 : boolean;
  signal type_cast_4316_inst_req_1 : boolean;
  signal phi_stmt_4132_req_1 : boolean;
  signal type_cast_4144_inst_req_0 : boolean;
  signal type_cast_4144_inst_ack_0 : boolean;
  signal type_cast_4144_inst_req_1 : boolean;
  signal type_cast_4144_inst_ack_1 : boolean;
  signal phi_stmt_4139_req_1 : boolean;
  signal type_cast_4150_inst_req_0 : boolean;
  signal type_cast_4150_inst_ack_0 : boolean;
  signal type_cast_4150_inst_req_1 : boolean;
  signal type_cast_4150_inst_ack_1 : boolean;
  signal phi_stmt_4145_req_1 : boolean;
  signal type_cast_4135_inst_req_0 : boolean;
  signal type_cast_4135_inst_ack_0 : boolean;
  signal type_cast_4135_inst_req_1 : boolean;
  signal type_cast_4135_inst_ack_1 : boolean;
  signal phi_stmt_4132_req_0 : boolean;
  signal type_cast_4701_inst_req_1 : boolean;
  signal type_cast_4701_inst_ack_1 : boolean;
  signal phi_stmt_4698_req_0 : boolean;
  signal type_cast_4694_inst_req_0 : boolean;
  signal type_cast_4694_inst_ack_0 : boolean;
  signal type_cast_4694_inst_req_1 : boolean;
  signal type_cast_4694_inst_ack_1 : boolean;
  signal phi_stmt_4691_req_0 : boolean;
  signal phi_stmt_4691_ack_0 : boolean;
  signal phi_stmt_4698_ack_0 : boolean;
  signal phi_stmt_4704_ack_0 : boolean;
  signal type_cast_4884_inst_req_0 : boolean;
  signal type_cast_4884_inst_ack_0 : boolean;
  signal type_cast_4884_inst_req_1 : boolean;
  signal type_cast_4884_inst_ack_1 : boolean;
  signal phi_stmt_4879_req_1 : boolean;
  signal type_cast_4876_inst_req_0 : boolean;
  signal type_cast_4876_inst_ack_0 : boolean;
  signal type_cast_4876_inst_req_1 : boolean;
  signal type_cast_4876_inst_ack_1 : boolean;
  signal phi_stmt_4873_req_0 : boolean;
  signal type_cast_4872_inst_req_0 : boolean;
  signal type_cast_4872_inst_ack_0 : boolean;
  signal type_cast_4872_inst_req_1 : boolean;
  signal type_cast_4872_inst_ack_1 : boolean;
  signal phi_stmt_4866_req_1 : boolean;
  signal type_cast_4882_inst_req_0 : boolean;
  signal type_cast_4882_inst_ack_0 : boolean;
  signal type_cast_4882_inst_req_1 : boolean;
  signal type_cast_4882_inst_ack_1 : boolean;
  signal phi_stmt_4879_req_0 : boolean;
  signal type_cast_4878_inst_req_0 : boolean;
  signal type_cast_4878_inst_ack_0 : boolean;
  signal type_cast_4878_inst_req_1 : boolean;
  signal type_cast_4878_inst_ack_1 : boolean;
  signal phi_stmt_4873_req_1 : boolean;
  signal phi_stmt_4866_req_0 : boolean;
  signal phi_stmt_4866_ack_0 : boolean;
  signal phi_stmt_4873_ack_0 : boolean;
  signal phi_stmt_4879_ack_0 : boolean;
  signal phi_stmt_5246_req_0 : boolean;
  signal type_cast_5258_inst_req_0 : boolean;
  signal type_cast_5258_inst_ack_0 : boolean;
  signal type_cast_5258_inst_req_1 : boolean;
  signal type_cast_5258_inst_ack_1 : boolean;
  signal phi_stmt_5253_req_1 : boolean;
  signal type_cast_5264_inst_req_0 : boolean;
  signal type_cast_5264_inst_ack_0 : boolean;
  signal type_cast_5264_inst_req_1 : boolean;
  signal type_cast_5264_inst_ack_1 : boolean;
  signal phi_stmt_5259_req_1 : boolean;
  signal type_cast_5252_inst_req_0 : boolean;
  signal type_cast_5252_inst_ack_0 : boolean;
  signal type_cast_5252_inst_req_1 : boolean;
  signal type_cast_5252_inst_ack_1 : boolean;
  signal phi_stmt_5246_req_1 : boolean;
  signal type_cast_5256_inst_req_0 : boolean;
  signal type_cast_5256_inst_ack_0 : boolean;
  signal type_cast_5256_inst_req_1 : boolean;
  signal type_cast_5256_inst_ack_1 : boolean;
  signal phi_stmt_5253_req_0 : boolean;
  signal type_cast_5262_inst_req_0 : boolean;
  signal type_cast_5262_inst_ack_0 : boolean;
  signal type_cast_5262_inst_req_1 : boolean;
  signal type_cast_5262_inst_ack_1 : boolean;
  signal phi_stmt_5259_req_0 : boolean;
  signal phi_stmt_5246_ack_0 : boolean;
  signal phi_stmt_5253_ack_0 : boolean;
  signal phi_stmt_5259_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_2152_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2152_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_2152_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_2152_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_2152: Block -- control-path 
    signal zeropad3D_CP_2152_elements: BooleanArray(1191 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_2152_elements(0) <= zeropad3D_CP_2152_start;
    zeropad3D_CP_2152_symbol <= zeropad3D_CP_2152_elements(819);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	16 
    -- CP-element group 0:  members (104) 
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773__entry__
      -- CP-element group 0: 	 branch_block_stmt_714/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/branch_block_stmt_714__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_update_start_
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/cr
      -- 
    crr_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => call_stmt_716_call_req_0); -- 
    ccr_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => call_stmt_716_call_req_1); -- 
    cr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => ptr_deref_727_load_0_req_1); -- 
    cr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => type_cast_731_inst_req_1); -- 
    cr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => STORE_row_high_733_store_0_req_1); -- 
    cr_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => ptr_deref_746_load_0_req_1); -- 
    cr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => type_cast_750_inst_req_1); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => STORE_col_high_752_store_0_req_1); -- 
    cr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => ptr_deref_765_load_0_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => type_cast_769_inst_req_1); -- 
    cr_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(0), ack => STORE_depth_high_771_store_0_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	863 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	824 
    -- CP-element group 1: 	825 
    -- CP-element group 1: 	827 
    -- CP-element group 1: 	828 
    -- CP-element group 1: 	830 
    -- CP-element group 1: 	831 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_714/merge_stmt_1306__exit__
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/cr
      -- 
    rr_11544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_905_inst_req_0); -- 
    cr_11549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_905_inst_req_1); -- 
    rr_11567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_912_inst_req_0); -- 
    cr_11572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_912_inst_req_1); -- 
    rr_11590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_919_inst_req_0); -- 
    cr_11595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1), ack => type_cast_919_inst_req_1); -- 
    zeropad3D_CP_2152_elements(1) <= zeropad3D_CP_2152_elements(863);
    -- CP-element group 2:  merge  fork  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	909 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	864 
    -- CP-element group 2: 	865 
    -- CP-element group 2: 	867 
    -- CP-element group 2: 	868 
    -- CP-element group 2: 	870 
    -- CP-element group 2: 	871 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_714/merge_stmt_1855__exit__
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Update/cr
      -- 
    rr_11867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1468_inst_req_0); -- 
    cr_11872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1468_inst_req_1); -- 
    rr_11890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1475_inst_req_0); -- 
    cr_11895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1475_inst_req_1); -- 
    rr_11913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1482_inst_req_0); -- 
    cr_11918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(2), ack => type_cast_1482_inst_req_1); -- 
    zeropad3D_CP_2152_elements(2) <= zeropad3D_CP_2152_elements(909);
    -- CP-element group 3:  merge  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	955 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	910 
    -- CP-element group 3: 	911 
    -- CP-element group 3: 	913 
    -- CP-element group 3: 	914 
    -- CP-element group 3: 	916 
    -- CP-element group 3: 	917 
    -- CP-element group 3:  members (27) 
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460
      -- CP-element group 3: 	 branch_block_stmt_714/merge_stmt_2420__exit__
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Update/cr
      -- 
    rr_12232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2018_inst_req_0); -- 
    cr_12237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2018_inst_req_1); -- 
    rr_12255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2031_inst_req_0); -- 
    cr_12260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2031_inst_req_1); -- 
    rr_12278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2027_inst_req_0); -- 
    cr_12283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(3), ack => type_cast_2027_inst_req_1); -- 
    zeropad3D_CP_2152_elements(3) <= zeropad3D_CP_2152_elements(955);
    -- CP-element group 4:  merge  fork  transition  place  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1003 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	956 
    -- CP-element group 4: 	957 
    -- CP-element group 4: 	959 
    -- CP-element group 4: 	960 
    -- CP-element group 4: 	962 
    -- CP-element group 4: 	963 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682
      -- CP-element group 4: 	 branch_block_stmt_714/merge_stmt_2981__exit__
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Update/cr
      -- 
    rr_12620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2602_inst_req_0); -- 
    rr_12597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2596_inst_req_0); -- 
    cr_12625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2602_inst_req_1); -- 
    cr_12602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2596_inst_req_1); -- 
    rr_12643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2608_inst_req_0); -- 
    cr_12648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(4), ack => type_cast_2608_inst_req_1); -- 
    zeropad3D_CP_2152_elements(4) <= zeropad3D_CP_2152_elements(1003);
    -- CP-element group 5:  merge  fork  transition  place  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1049 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	1004 
    -- CP-element group 5: 	1005 
    -- CP-element group 5: 	1007 
    -- CP-element group 5: 	1008 
    -- CP-element group 5: 	1010 
    -- CP-element group 5: 	1011 
    -- CP-element group 5:  members (27) 
      -- CP-element group 5: 	 branch_block_stmt_714/merge_stmt_3558__exit__
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Update/cr
      -- 
    rr_12977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3157_inst_req_0); -- 
    cr_12982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3157_inst_req_1); -- 
    rr_13000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3153_inst_req_0); -- 
    cr_13005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3153_inst_req_1); -- 
    rr_13023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3144_inst_req_0); -- 
    cr_13028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(5), ack => type_cast_3144_inst_req_1); -- 
    zeropad3D_CP_2152_elements(5) <= zeropad3D_CP_2152_elements(1049);
    -- CP-element group 6:  merge  fork  transition  place  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1097 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	1050 
    -- CP-element group 6: 	1051 
    -- CP-element group 6: 	1053 
    -- CP-element group 6: 	1054 
    -- CP-element group 6: 	1056 
    -- CP-element group 6: 	1057 
    -- CP-element group 6:  members (27) 
      -- CP-element group 6: 	 branch_block_stmt_714/merge_stmt_4131__exit__
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Update/cr
      -- 
    rr_13342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3731_inst_req_0); -- 
    cr_13347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3731_inst_req_1); -- 
    rr_13365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3740_inst_req_0); -- 
    cr_13370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3740_inst_req_1); -- 
    rr_13388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3744_inst_req_0); -- 
    cr_13393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(6), ack => type_cast_3744_inst_req_1); -- 
    zeropad3D_CP_2152_elements(6) <= zeropad3D_CP_2152_elements(1097);
    -- CP-element group 7:  merge  fork  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1143 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	1098 
    -- CP-element group 7: 	1099 
    -- CP-element group 7: 	1101 
    -- CP-element group 7: 	1102 
    -- CP-element group 7: 	1104 
    -- CP-element group 7: 	1105 
    -- CP-element group 7:  members (27) 
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341
      -- CP-element group 7: 	 branch_block_stmt_714/merge_stmt_4690__exit__
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Update/cr
      -- 
    rr_13722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4303_inst_req_0); -- 
    cr_13727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4303_inst_req_1); -- 
    rr_13768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4316_inst_req_0); -- 
    cr_13750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4309_inst_req_1); -- 
    rr_13745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4309_inst_req_0); -- 
    cr_13773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(7), ack => type_cast_4316_inst_req_1); -- 
    zeropad3D_CP_2152_elements(7) <= zeropad3D_CP_2152_elements(1143);
    -- CP-element group 8:  merge  fork  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1191 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	1144 
    -- CP-element group 8: 	1145 
    -- CP-element group 8: 	1147 
    -- CP-element group 8: 	1148 
    -- CP-element group 8: 	1150 
    -- CP-element group 8: 	1151 
    -- CP-element group 8:  members (27) 
      -- CP-element group 8: 	 branch_block_stmt_714/merge_stmt_5245__exit__
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Update/cr
      -- 
    rr_14087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4884_inst_req_0); -- 
    cr_14092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4884_inst_req_1); -- 
    rr_14110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4876_inst_req_0); -- 
    cr_14115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4876_inst_req_1); -- 
    rr_14133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4872_inst_req_0); -- 
    cr_14138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(8), ack => type_cast_4872_inst_req_1); -- 
    zeropad3D_CP_2152_elements(8) <= zeropad3D_CP_2152_elements(1191);
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Sample/cra
      -- 
    cra_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_716_call_ack_0, ack => zeropad3D_CP_2152_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	36 
    -- CP-element group 10: 	37 
    -- CP-element group 10: 	38 
    -- CP-element group 10: 	39 
    -- CP-element group 10: 	40 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_Update/cca
      -- 
    cca_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_716_call_ack_1, ack => zeropad3D_CP_2152_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/$entry
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/$entry
      -- CP-element group 11: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/rr
      -- 
    rr_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(11), ack => ptr_deref_727_load_0_req_0); -- 
    zeropad3D_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(37) & zeropad3D_CP_2152_elements(0);
      gj_zeropad3D_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/$exit
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Sample/word_access_start/word_0/ra
      -- 
    ra_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_727_load_0_ack_0, ack => zeropad3D_CP_2152_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/$entry
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/$exit
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/merge_req
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_727_Update/ptr_deref_727_Merge/merge_ack
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/rr
      -- 
    ca_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_727_load_0_ack_1, ack => zeropad3D_CP_2152_elements(13)); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(13), ack => type_cast_731_inst_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Sample/ra
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_0, ack => zeropad3D_CP_2152_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_731_Update/ca
      -- 
    ca_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_731_inst_ack_1, ack => zeropad3D_CP_2152_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	40 
    -- CP-element group 16: 	15 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/$exit
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/split_req
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/STORE_row_high_733_Split/split_ack
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/rr
      -- 
    rr_2699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(16), ack => STORE_row_high_733_store_0_req_0); -- 
    zeropad3D_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(40) & zeropad3D_CP_2152_elements(15) & zeropad3D_CP_2152_elements(0);
      gj_zeropad3D_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Sample/word_access_start/word_0/ra
      -- 
    ra_2700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_733_store_0_ack_0, ack => zeropad3D_CP_2152_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_row_high_733_Update/word_access_complete/word_0/ca
      -- 
    ca_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_row_high_733_store_0_ack_1, ack => zeropad3D_CP_2152_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	38 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/rr
      -- 
    rr_2744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(19), ack => ptr_deref_746_load_0_req_0); -- 
    zeropad3D_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(38) & zeropad3D_CP_2152_elements(0);
      gj_zeropad3D_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Sample/word_access_start/word_0/ra
      -- 
    ra_2745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_746_load_0_ack_0, ack => zeropad3D_CP_2152_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (12) 
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/$entry
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/$exit
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/merge_req
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_746_Update/ptr_deref_746_Merge/merge_ack
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/rr
      -- 
    ca_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_746_load_0_ack_1, ack => zeropad3D_CP_2152_elements(21)); -- 
    rr_2769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(21), ack => type_cast_750_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Sample/ra
      -- 
    ra_2770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => zeropad3D_CP_2152_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_750_Update/ca
      -- 
    ca_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => zeropad3D_CP_2152_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	35 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/$exit
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/split_req
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/STORE_col_high_752_Split/split_ack
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/$entry
      -- CP-element group 24: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/rr
      -- 
    rr_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(24), ack => STORE_col_high_752_store_0_req_0); -- 
    zeropad3D_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(23) & zeropad3D_CP_2152_elements(35) & zeropad3D_CP_2152_elements(0);
      gj_zeropad3D_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Sample/word_access_start/word_0/ra
      -- 
    ra_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_752_store_0_ack_0, ack => zeropad3D_CP_2152_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	41 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_col_high_752_Update/word_access_complete/word_0/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_col_high_752_store_0_ack_1, ack => zeropad3D_CP_2152_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	39 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/$entry
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/$entry
      -- CP-element group 27: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/rr
      -- 
    rr_2841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(27), ack => ptr_deref_765_load_0_req_0); -- 
    zeropad3D_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(39) & zeropad3D_CP_2152_elements(0);
      gj_zeropad3D_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/$exit
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Sample/word_access_start/word_0/ra
      -- 
    ra_2842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_765_load_0_ack_0, ack => zeropad3D_CP_2152_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (12) 
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/word_access_complete/word_0/ca
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/$entry
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/$exit
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/merge_req
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/ptr_deref_765_Update/ptr_deref_765_Merge/merge_ack
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/rr
      -- 
    ca_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_765_load_0_ack_1, ack => zeropad3D_CP_2152_elements(29)); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(29), ack => type_cast_769_inst_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_0, ack => zeropad3D_CP_2152_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/type_cast_769_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_769_inst_ack_1, ack => zeropad3D_CP_2152_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	36 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/$exit
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/split_req
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/STORE_depth_high_771_Split/split_ack
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/rr
      -- 
    rr_2893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(32), ack => STORE_depth_high_771_store_0_req_0); -- 
    zeropad3D_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(31) & zeropad3D_CP_2152_elements(36) & zeropad3D_CP_2152_elements(0);
      gj_zeropad3D_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Sample/word_access_start/word_0/ra
      -- 
    ra_2894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_771_store_0_ack_0, ack => zeropad3D_CP_2152_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/STORE_depth_high_771_Update/word_access_complete/word_0/ca
      -- 
    ca_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_depth_high_771_store_0_ack_1, ack => zeropad3D_CP_2152_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	24 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_STORE_col_high_752_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  transition  delay-element  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	10 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	32 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_STORE_depth_high_771_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(36) is a control-delay.
    cp_element_36_delay: control_delay_element  generic map(name => " 36_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(36), clk => clk, reset =>reset);
    -- CP-element group 37:  transition  delay-element  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	10 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_ptr_deref_727_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(37) is a control-delay.
    cp_element_37_delay: control_delay_element  generic map(name => " 37_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(37), clk => clk, reset =>reset);
    -- CP-element group 38:  transition  delay-element  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	10 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	19 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_ptr_deref_746_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(38) is a control-delay.
    cp_element_38_delay: control_delay_element  generic map(name => " 38_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(38), clk => clk, reset =>reset);
    -- CP-element group 39:  transition  delay-element  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	10 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	27 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_ptr_deref_765_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(39) is a control-delay.
    cp_element_39_delay: control_delay_element  generic map(name => " 39_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(39), clk => clk, reset =>reset);
    -- CP-element group 40:  transition  delay-element  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	16 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/call_stmt_716_STORE_row_high_733_delay
      -- 
    -- Element group zeropad3D_CP_2152_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(10), ack => zeropad3D_CP_2152_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: 	26 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	44 
    -- CP-element group 41: 	45 
    -- CP-element group 41: 	46 
    -- CP-element group 41: 	47 
    -- CP-element group 41: 	48 
    -- CP-element group 41: 	49 
    -- CP-element group 41: 	50 
    -- CP-element group 41: 	51 
    -- CP-element group 41: 	53 
    -- CP-element group 41: 	55 
    -- CP-element group 41: 	57 
    -- CP-element group 41:  members (101) 
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896__entry__
      -- CP-element group 41: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773__exit__
      -- CP-element group 41: 	 branch_block_stmt_714/call_stmt_716_to_assign_stmt_773/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_update_start_
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/cr
      -- 
    rr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_pad_776_load_0_req_0); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_pad_776_load_0_req_1); -- 
    rr_2963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_depth_high_779_load_0_req_0); -- 
    cr_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_depth_high_779_load_0_req_1); -- 
    rr_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_col_high_782_load_0_req_0); -- 
    cr_3007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => LOAD_col_high_782_load_0_req_1); -- 
    rr_3046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_794_load_0_req_0); -- 
    cr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_794_load_0_req_1); -- 
    rr_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_806_load_0_req_0); -- 
    cr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => ptr_deref_806_load_0_req_1); -- 
    cr_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => type_cast_810_inst_req_1); -- 
    cr_3140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => type_cast_814_inst_req_1); -- 
    cr_3154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(41), ack => type_cast_854_inst_req_1); -- 
    zeropad3D_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(18) & zeropad3D_CP_2152_elements(26) & zeropad3D_CP_2152_elements(34);
      gj_zeropad3D_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Sample/word_access_start/word_0/ra
      -- 
    ra_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_776_load_0_ack_0, ack => zeropad3D_CP_2152_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/$entry
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/$exit
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/merge_req
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_pad_776_Update/LOAD_pad_776_Merge/merge_ack
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/rr
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_776_load_0_ack_1, ack => zeropad3D_CP_2152_elements(43)); -- 
    rr_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(43), ack => type_cast_854_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	41 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/$exit
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Sample/word_access_start/word_0/ra
      -- 
    ra_2964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_779_load_0_ack_0, ack => zeropad3D_CP_2152_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	41 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	52 
    -- CP-element group 45:  members (12) 
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/word_access_complete/word_0/ca
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/$entry
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/$exit
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/merge_req
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_depth_high_779_Update/LOAD_depth_high_779_Merge/merge_ack
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/rr
      -- 
    ca_2975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_779_load_0_ack_1, ack => zeropad3D_CP_2152_elements(45)); -- 
    rr_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(45), ack => type_cast_810_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	41 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/$exit
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Sample/word_access_start/word_0/ra
      -- 
    ra_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_782_load_0_ack_0, ack => zeropad3D_CP_2152_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	41 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	54 
    -- CP-element group 47:  members (12) 
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/$entry
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/$exit
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/merge_req
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/LOAD_col_high_782_Update/LOAD_col_high_782_Merge/merge_ack
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/rr
      -- 
    ca_3008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_782_load_0_ack_1, ack => zeropad3D_CP_2152_elements(47)); -- 
    rr_3135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(47), ack => type_cast_814_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	41 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/$exit
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Sample/word_access_start/word_0/ra
      -- 
    ra_3047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_794_load_0_ack_0, ack => zeropad3D_CP_2152_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	41 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/word_access_complete/word_0/ca
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/$entry
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/$exit
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/merge_req
      -- CP-element group 49: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_794_Update/ptr_deref_794_Merge/merge_ack
      -- 
    ca_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_794_load_0_ack_1, ack => zeropad3D_CP_2152_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Sample/word_access_start/word_0/ra
      -- 
    ra_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_806_load_0_ack_0, ack => zeropad3D_CP_2152_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	41 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	58 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/$entry
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/$exit
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/merge_req
      -- CP-element group 51: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/ptr_deref_806_Update/ptr_deref_806_Merge/merge_ack
      -- 
    ca_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_806_load_0_ack_1, ack => zeropad3D_CP_2152_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	45 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Sample/ra
      -- 
    ra_3122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_810_inst_ack_0, ack => zeropad3D_CP_2152_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	41 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	58 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_810_Update/ca
      -- 
    ca_3127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_810_inst_ack_1, ack => zeropad3D_CP_2152_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	47 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Sample/ra
      -- 
    ra_3136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_0, ack => zeropad3D_CP_2152_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	41 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_814_Update/ca
      -- 
    ca_3141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_1, ack => zeropad3D_CP_2152_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Sample/ra
      -- 
    ra_3150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => zeropad3D_CP_2152_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/type_cast_854_Update/ca
      -- 
    ca_3155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => zeropad3D_CP_2152_elements(57)); -- 
    -- CP-element group 58:  join  fork  transition  place  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	51 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	820 
    -- CP-element group 58: 	821 
    -- CP-element group 58: 	822 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody
      -- CP-element group 58: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896__exit__
      -- CP-element group 58: 	 branch_block_stmt_714/assign_stmt_777_to_assign_stmt_896/$exit
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/$entry
      -- CP-element group 58: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$entry
      -- 
    zeropad3D_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(49) & zeropad3D_CP_2152_elements(51) & zeropad3D_CP_2152_elements(53) & zeropad3D_CP_2152_elements(55) & zeropad3D_CP_2152_elements(57);
      gj_zeropad3D_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	838 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/ra
      -- 
    ra_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_0, ack => zeropad3D_CP_2152_elements(59)); -- 
    -- CP-element group 60:  branch  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	838 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933__entry__
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932__exit__
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/$exit
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_714/R_cmp_934_place
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_714/if_stmt_933_else_link/$entry
      -- 
    ca_3172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_924_inst_ack_1, ack => zeropad3D_CP_2152_elements(60)); -- 
    branch_req_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(60), ack => if_stmt_933_branch_req_0); -- 
    -- CP-element group 61:  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	839 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_714/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_714/if_stmt_933_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_714/if_stmt_933_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_714/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_714/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_933_branch_ack_1, ack => zeropad3D_CP_2152_elements(61)); -- 
    -- CP-element group 62:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	66 
    -- CP-element group 62:  members (27) 
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939__exit__
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964__entry__
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_update_start_
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_update_start_
      -- CP-element group 62: 	 branch_block_stmt_714/whilex_xbody_lorx_xlhsx_xfalse
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/rr
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/cr
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/if_stmt_933_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_714/if_stmt_933_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_714/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/whilex_xbody_lorx_xlhsx_xfalse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_714/merge_stmt_939_PhiAck/dummy
      -- 
    else_choice_transition_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_933_branch_ack_0, ack => zeropad3D_CP_2152_elements(62)); -- 
    rr_3210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(62), ack => LOAD_row_high_941_load_0_req_0); -- 
    cr_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(62), ack => LOAD_row_high_941_load_0_req_1); -- 
    cr_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(62), ack => type_cast_945_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/ra
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Sample/word_access_start/$exit
      -- 
    ra_3211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_941_load_0_ack_0, ack => zeropad3D_CP_2152_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (12) 
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/merge_ack
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/LOAD_row_high_941_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/LOAD_row_high_941_Update/word_access_complete/word_0/$exit
      -- 
    ca_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_941_load_0_ack_1, ack => zeropad3D_CP_2152_elements(64)); -- 
    rr_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(64), ack => type_cast_945_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Sample/ra
      -- 
    ra_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_0, ack => zeropad3D_CP_2152_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964__exit__
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965__entry__
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_714/R_cmp56_966_place
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/$exit
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/if_stmt_965_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_714/assign_stmt_942_to_assign_stmt_964/type_cast_945_Update/$exit
      -- 
    ca_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_945_inst_ack_1, ack => zeropad3D_CP_2152_elements(66)); -- 
    branch_req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(66), ack => if_stmt_965_branch_req_0); -- 
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (18) 
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971__exit__
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983__entry__
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse58
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_update_start_
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_714/if_stmt_965_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_714/if_stmt_965_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse58_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_lorx_xlhsx_xfalse58_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_714/merge_stmt_971_PhiAck/dummy
      -- 
    if_choice_transition_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_965_branch_ack_1, ack => zeropad3D_CP_2152_elements(67)); -- 
    cr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(67), ack => type_cast_975_inst_req_1); -- 
    rr_3271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(67), ack => type_cast_975_inst_req_0); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	839 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_ifx_xthen
      -- CP-element group 68: 	 branch_block_stmt_714/if_stmt_965_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_714/if_stmt_965_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_714/lorx_xlhsx_xfalse_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_965_branch_ack_0, ack => zeropad3D_CP_2152_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_sample_completed_
      -- 
    ra_3272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_0, ack => zeropad3D_CP_2152_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_714/R_cmp63_985_place
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983__exit__
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984__entry__
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/type_cast_975_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_714/assign_stmt_976_to_assign_stmt_983/$exit
      -- CP-element group 70: 	 branch_block_stmt_714/if_stmt_984_else_link/$entry
      -- 
    ca_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_1, ack => zeropad3D_CP_2152_elements(70)); -- 
    branch_req_3285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(70), ack => if_stmt_984_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	839 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_714/if_stmt_984_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_714/if_stmt_984_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_ifx_xthen
      -- CP-element group 71: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_ifx_xthen_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_ifx_xthen_PhiReq/$exit
      -- 
    if_choice_transition_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_984_branch_ack_1, ack => zeropad3D_CP_2152_elements(71)); -- 
    -- CP-element group 72:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	76 
    -- CP-element group 72:  members (27) 
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015__entry__
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990__exit__
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_update_start_
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/cr
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/rr
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_update_start_
      -- CP-element group 72: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_lorx_xlhsx_xfalse65
      -- CP-element group 72: 	 branch_block_stmt_714/if_stmt_984_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_714/if_stmt_984_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_lorx_xlhsx_xfalse65_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/lorx_xlhsx_xfalse58_lorx_xlhsx_xfalse65_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_714/merge_stmt_990_PhiAck/dummy
      -- 
    else_choice_transition_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_984_branch_ack_0, ack => zeropad3D_CP_2152_elements(72)); -- 
    cr_3345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(72), ack => type_cast_996_inst_req_1); -- 
    cr_3326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(72), ack => LOAD_col_high_992_load_0_req_1); -- 
    rr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(72), ack => LOAD_col_high_992_load_0_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/ra
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/word_access_start/$exit
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_sample_completed_
      -- 
    ra_3316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_992_load_0_ack_0, ack => zeropad3D_CP_2152_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (12) 
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/merge_ack
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/merge_req
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/LOAD_col_high_992_Merge/$entry
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/ca
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/word_access_complete/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/LOAD_col_high_992_update_completed_
      -- 
    ca_3327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_992_load_0_ack_1, ack => zeropad3D_CP_2152_elements(74)); -- 
    rr_3340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(74), ack => type_cast_996_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_sample_completed_
      -- 
    ra_3341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_0, ack => zeropad3D_CP_2152_elements(75)); -- 
    -- CP-element group 76:  branch  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	72 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (13) 
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016__entry__
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015__exit__
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_else_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_if_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/R_cmp74_1017_place
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_eval_test/branch_req
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_eval_test/$exit
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_eval_test/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/if_stmt_1016_dead_link/$entry
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/type_cast_996_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_714/assign_stmt_993_to_assign_stmt_1015/$exit
      -- 
    ca_3346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_1, ack => zeropad3D_CP_2152_elements(76)); -- 
    branch_req_3354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(76), ack => if_stmt_1016_branch_req_0); -- 
    -- CP-element group 77:  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	93 
    -- CP-element group 77: 	94 
    -- CP-element group 77: 	96 
    -- CP-element group 77: 	98 
    -- CP-element group 77: 	100 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	104 
    -- CP-element group 77: 	106 
    -- CP-element group 77: 	108 
    -- CP-element group 77: 	111 
    -- CP-element group 77:  members (46) 
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186__entry__
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081__exit__
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xelse
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/if_stmt_1016_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/if_stmt_1016_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/req
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_update_start_
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xelse_PhiReq/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xelse_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_714/merge_stmt_1081_PhiAck/dummy
      -- 
    if_choice_transition_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1016_branch_ack_1, ack => zeropad3D_CP_2152_elements(77)); -- 
    cr_3536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1149_inst_req_1); -- 
    req_3582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => addr_of_1156_final_reg_req_1); -- 
    cr_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => ptr_deref_1160_load_0_req_1); -- 
    cr_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1085_inst_req_1); -- 
    cr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1174_inst_req_1); -- 
    rr_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => type_cast_1085_inst_req_0); -- 
    req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => array_obj_ref_1155_index_offset_req_1); -- 
    req_3677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => array_obj_ref_1180_index_offset_req_1); -- 
    req_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => addr_of_1181_final_reg_req_1); -- 
    cr_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(77), ack => ptr_deref_1184_store_0_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	839 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xthen
      -- CP-element group 78: 	 branch_block_stmt_714/if_stmt_1016_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_714/if_stmt_1016_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xthen_PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_714/lorx_xlhsx_xfalse65_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1016_branch_ack_0, ack => zeropad3D_CP_2152_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	839 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/$exit
      -- 
    ra_3377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1026_inst_ack_0, ack => zeropad3D_CP_2152_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	839 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/$exit
      -- 
    ca_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1026_inst_ack_1, ack => zeropad3D_CP_2152_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	839 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_sample_completed_
      -- 
    ra_3391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1031_inst_ack_0, ack => zeropad3D_CP_2152_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	839 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/$exit
      -- 
    ca_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1031_inst_ack_1, ack => zeropad3D_CP_2152_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_sample_start_
      -- 
    rr_3404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(83), ack => type_cast_1066_inst_req_0); -- 
    zeropad3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(80) & zeropad3D_CP_2152_elements(82);
      gj_zeropad3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_sample_completed_
      -- 
    ra_3405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_0, ack => zeropad3D_CP_2152_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	839 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (16) 
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/scale_rename_ack
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/scale_rename_req
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/$exit
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scale_1/$entry
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/index_resize_ack
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/index_resize_req
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/$exit
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resize_1/$entry
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_computed_1
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_scaled_1
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_index_resized_1
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/$entry
      -- 
    ca_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_1, ack => zeropad3D_CP_2152_elements(85)); -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(85), ack => array_obj_ref_1072_index_offset_req_0); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	92 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_sample_complete
      -- CP-element group 86: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Sample/$exit
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1072_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	839 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (11) 
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_offset_calculated
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_root_address_calculated
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/req
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/$entry
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/sum_rename_ack
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/sum_rename_req
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/$exit
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_base_plus_offset/$entry
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/ack
      -- CP-element group 87: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/$exit
      -- 
    ack_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1072_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(87)); -- 
    req_3450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(87), ack => addr_of_1073_final_reg_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/ack
      -- CP-element group 88: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_request/$exit
      -- 
    ack_3451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1073_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	839 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (28) 
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/split_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/ptr_deref_1076_Split/split_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/root_register_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/root_register_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_addrgen/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/sum_rename_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/sum_rename_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_plus_offset/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/base_resize_ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/base_resize_req
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_addr_resize/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_address_resized
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_root_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_word_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_base_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/rr
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/ack
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/$entry
      -- 
    ack_3456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1073_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(89)); -- 
    rr_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(89), ack => ptr_deref_1076_store_0_req_0); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/$exit
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/ra
      -- CP-element group 90: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Sample/word_access_start/word_0/$exit
      -- 
    ra_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_store_0_ack_0, ack => zeropad3D_CP_2152_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	839 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/$exit
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/ca
      -- 
    ca_3506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_store_0_ack_1, ack => zeropad3D_CP_2152_elements(91)); -- 
    -- CP-element group 92:  join  transition  place  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	86 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	840 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079__exit__
      -- CP-element group 92: 	 branch_block_stmt_714/ifx_xthen_ifx_xend
      -- CP-element group 92: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/$exit
      -- CP-element group 92: 	 branch_block_stmt_714/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 92: 	 branch_block_stmt_714/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(86) & zeropad3D_CP_2152_elements(91);
      gj_zeropad3D_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	77 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_sample_completed_
      -- 
    ra_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_0, ack => zeropad3D_CP_2152_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	77 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	103 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1085_update_completed_
      -- 
    ca_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1085_inst_ack_1, ack => zeropad3D_CP_2152_elements(94)); -- 
    rr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(94), ack => type_cast_1149_inst_req_0); -- 
    rr_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(94), ack => type_cast_1174_inst_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_sample_completed_
      -- 
    ra_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_0, ack => zeropad3D_CP_2152_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	77 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (16) 
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/scale_rename_ack
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/scale_rename_req
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1149_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/$exit
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scale_1/$entry
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/index_resize_ack
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/index_resize_req
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/$exit
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resize_1/$entry
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_computed_1
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_scaled_1
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_index_resized_1
      -- CP-element group 96: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/req
      -- 
    ca_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_1, ack => zeropad3D_CP_2152_elements(96)); -- 
    req_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(96), ack => array_obj_ref_1155_index_offset_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	112 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_sample_complete
      -- CP-element group 97: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Sample/ack
      -- 
    ack_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1155_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	77 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (11) 
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/req
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_offset_calculated
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_root_address_calculated
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/$entry
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/sum_rename_ack
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/sum_rename_req
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/$exit
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_base_plus_offset/$entry
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/ack
      -- CP-element group 98: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1155_final_index_sum_regn_Update/$exit
      -- 
    ack_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1155_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(98)); -- 
    req_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(98), ack => addr_of_1156_final_reg_req_0); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/ack
      -- CP-element group 99: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_request/$exit
      -- CP-element group 99: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_sample_completed_
      -- 
    ack_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1156_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	77 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (24) 
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_root_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/root_register_ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/root_register_req
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_word_addrgen/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/sum_rename_ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/sum_rename_req
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_plus_offset/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/base_resize_ack
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/base_resize_req
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/$exit
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_addr_resize/$entry
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1156_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_base_address_resized
      -- CP-element group 100: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/rr
      -- 
    ack_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1156_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(100)); -- 
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(100), ack => ptr_deref_1160_load_0_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Sample/word_access_start/$exit
      -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1160_load_0_ack_0, ack => zeropad3D_CP_2152_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	109 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/ptr_deref_1160_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1160_Update/word_access_complete/word_0/$exit
      -- 
    ca_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1160_load_0_ack_1, ack => zeropad3D_CP_2152_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	94 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Sample/$exit
      -- 
    ra_3642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_0, ack => zeropad3D_CP_2152_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	77 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (16) 
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/type_cast_1174_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resized_1
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scaled_1
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_computed_1
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/$entry
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/$exit
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/index_resize_req
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_resize_1/index_resize_ack
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/$entry
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/$exit
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/scale_rename_req
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_index_scale_1/scale_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/req
      -- 
    ca_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_1, ack => zeropad3D_CP_2152_elements(104)); -- 
    req_3672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(104), ack => array_obj_ref_1180_index_offset_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_sample_complete
      -- CP-element group 105: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Sample/ack
      -- 
    ack_3673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1180_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	77 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (11) 
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/$entry
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_root_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_offset_calculated
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_final_index_sum_regn_Update/ack
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/$entry
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/$exit
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/sum_rename_req
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/array_obj_ref_1180_base_plus_offset/sum_rename_ack
      -- CP-element group 106: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/req
      -- 
    ack_3678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1180_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(106)); -- 
    req_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(106), ack => addr_of_1181_final_reg_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/$exit
      -- CP-element group 107: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_request/ack
      -- 
    ack_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1181_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(107)); -- 
    -- CP-element group 108:  fork  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	77 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (19) 
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/addr_of_1181_complete/ack
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_root_address_calculated
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_address_resized
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/$entry
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/base_resize_req
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_addr_resize/base_resize_ack
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/$entry
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/sum_rename_req
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_base_plus_offset/sum_rename_ack
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/$entry
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/$exit
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/root_register_req
      -- CP-element group 108: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_word_addrgen/root_register_ack
      -- 
    ack_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1181_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	102 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/$exit
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/split_req
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/ptr_deref_1184_Split/split_ack
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/$entry
      -- CP-element group 109: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/rr
      -- 
    rr_3731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(109), ack => ptr_deref_1184_store_0_req_0); -- 
    zeropad3D_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(102) & zeropad3D_CP_2152_elements(108);
      gj_zeropad3D_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Sample/word_access_start/word_0/ra
      -- 
    ra_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1184_store_0_ack_0, ack => zeropad3D_CP_2152_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	77 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/ptr_deref_1184_Update/word_access_complete/word_0/ca
      -- 
    ca_3743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1184_store_0_ack_1, ack => zeropad3D_CP_2152_elements(111)); -- 
    -- CP-element group 112:  join  transition  place  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	97 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	840 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_714/ifx_xelse_ifx_xend
      -- CP-element group 112: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186__exit__
      -- CP-element group 112: 	 branch_block_stmt_714/assign_stmt_1086_to_assign_stmt_1186/$exit
      -- CP-element group 112: 	 branch_block_stmt_714/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 112: 	 branch_block_stmt_714/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(97) & zeropad3D_CP_2152_elements(105) & zeropad3D_CP_2152_elements(111);
      gj_zeropad3D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	840 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/ra
      -- 
    ra_3755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_0, ack => zeropad3D_CP_2152_elements(113)); -- 
    -- CP-element group 114:  branch  transition  place  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	840 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (13) 
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207__entry__
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206__exit__
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/$exit
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_dead_link/$entry
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_eval_test/$entry
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_eval_test/$exit
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_eval_test/branch_req
      -- CP-element group 114: 	 branch_block_stmt_714/R_cmp143_1208_place
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_if_link/$entry
      -- CP-element group 114: 	 branch_block_stmt_714/if_stmt_1207_else_link/$entry
      -- 
    ca_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_1, ack => zeropad3D_CP_2152_elements(114)); -- 
    branch_req_3768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(114), ack => if_stmt_1207_branch_req_0); -- 
    -- CP-element group 115:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	849 
    -- CP-element group 115: 	850 
    -- CP-element group 115: 	852 
    -- CP-element group 115: 	853 
    -- CP-element group 115: 	855 
    -- CP-element group 115: 	856 
    -- CP-element group 115:  members (40) 
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219__entry__
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213__exit__
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219__exit__
      -- CP-element group 115: 	 branch_block_stmt_714/if_stmt_1207_if_link/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/if_stmt_1207_if_link/if_choice_transition
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xend_ifx_xthen145
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/assign_stmt_1219/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xend_ifx_xthen145_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xend_ifx_xthen145_PhiReq/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_714/merge_stmt_1213_PhiAck/dummy
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/cr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/cr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1207_branch_ack_1, ack => zeropad3D_CP_2152_elements(115)); -- 
    rr_11780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1316_inst_req_0); -- 
    cr_11785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1316_inst_req_1); -- 
    rr_11803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1325_inst_req_0); -- 
    cr_11808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1325_inst_req_1); -- 
    rr_11826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1312_inst_req_0); -- 
    cr_11831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(115), ack => type_cast_1312_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  place  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116: 	119 
    -- CP-element group 116: 	120 
    -- CP-element group 116: 	122 
    -- CP-element group 116: 	125 
    -- CP-element group 116: 	127 
    -- CP-element group 116: 	128 
    -- CP-element group 116: 	129 
    -- CP-element group 116: 	131 
    -- CP-element group 116:  members (54) 
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221__exit__
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299__entry__
      -- CP-element group 116: 	 branch_block_stmt_714/if_stmt_1207_else_link/$exit
      -- CP-element group 116: 	 branch_block_stmt_714/if_stmt_1207_else_link/else_choice_transition
      -- CP-element group 116: 	 branch_block_stmt_714/ifx_xend_ifx_xelse150
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/cr
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_update_start_
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_714/ifx_xend_ifx_xelse150_PhiReq/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/ifx_xend_ifx_xelse150_PhiReq/$exit
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiReqMerge
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiAck/$entry
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiAck/$exit
      -- CP-element group 116: 	 branch_block_stmt_714/merge_stmt_1221_PhiAck/dummy
      -- 
    else_choice_transition_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1207_branch_ack_0, ack => zeropad3D_CP_2152_elements(116)); -- 
    rr_3793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1231_inst_req_0); -- 
    cr_3798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1231_inst_req_1); -- 
    rr_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_col_high_1234_load_0_req_0); -- 
    cr_3826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_col_high_1234_load_0_req_1); -- 
    cr_3845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1238_inst_req_1); -- 
    cr_3859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1258_inst_req_1); -- 
    cr_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1275_inst_req_1); -- 
    rr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_row_high_1278_load_0_req_0); -- 
    cr_3901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => LOAD_row_high_1278_load_0_req_1); -- 
    cr_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(116), ack => type_cast_1282_inst_req_1); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Sample/ra
      -- 
    ra_3794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => zeropad3D_CP_2152_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1231_Update/ca
      -- 
    ca_3799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => zeropad3D_CP_2152_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Sample/word_access_start/word_0/ra
      -- 
    ra_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1234_load_0_ack_0, ack => zeropad3D_CP_2152_elements(119)); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	116 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (12) 
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_col_high_1234_Update/LOAD_col_high_1234_Merge/merge_ack
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/rr
      -- 
    ca_3827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1234_load_0_ack_1, ack => zeropad3D_CP_2152_elements(120)); -- 
    rr_3840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(120), ack => type_cast_1238_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Sample/ra
      -- 
    ra_3841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => zeropad3D_CP_2152_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	116 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1238_Update/ca
      -- 
    ca_3846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => zeropad3D_CP_2152_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/rr
      -- 
    rr_3854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(123), ack => type_cast_1258_inst_req_0); -- 
    zeropad3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(118) & zeropad3D_CP_2152_elements(122);
      gj_zeropad3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Sample/ra
      -- 
    ra_3855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_0, ack => zeropad3D_CP_2152_elements(124)); -- 
    -- CP-element group 125:  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	116 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (6) 
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1258_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/rr
      -- 
    ca_3860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_1, ack => zeropad3D_CP_2152_elements(125)); -- 
    rr_3868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(125), ack => type_cast_1275_inst_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Sample/ra
      -- 
    ra_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_0, ack => zeropad3D_CP_2152_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	116 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	132 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1275_Update/ca
      -- 
    ca_3874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_1, ack => zeropad3D_CP_2152_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	116 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/$exit
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/$exit
      -- CP-element group 128: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Sample/word_access_start/word_0/ra
      -- 
    ra_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1278_load_0_ack_0, ack => zeropad3D_CP_2152_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	116 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (12) 
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/word_access_complete/word_0/ca
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/$entry
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/$exit
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/merge_req
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/LOAD_row_high_1278_Update/LOAD_row_high_1278_Merge/merge_ack
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/rr
      -- 
    ca_3902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1278_load_0_ack_1, ack => zeropad3D_CP_2152_elements(129)); -- 
    rr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(129), ack => type_cast_1282_inst_req_0); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Sample/ra
      -- 
    ra_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1282_inst_ack_0, ack => zeropad3D_CP_2152_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	116 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/type_cast_1282_Update/ca
      -- 
    ca_3921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1282_inst_ack_1, ack => zeropad3D_CP_2152_elements(131)); -- 
    -- CP-element group 132:  branch  join  transition  place  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	127 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (10) 
      -- CP-element group 132: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299__exit__
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300__entry__
      -- CP-element group 132: 	 branch_block_stmt_714/assign_stmt_1227_to_assign_stmt_1299/$exit
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_dead_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_eval_test/$entry
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_eval_test/$exit
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_eval_test/branch_req
      -- CP-element group 132: 	 branch_block_stmt_714/R_cmp176_1301_place
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_if_link/$entry
      -- CP-element group 132: 	 branch_block_stmt_714/if_stmt_1300_else_link/$entry
      -- 
    branch_req_3929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(132), ack => if_stmt_1300_branch_req_0); -- 
    zeropad3D_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(127) & zeropad3D_CP_2152_elements(131);
      gj_zeropad3D_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	136 
    -- CP-element group 133: 	138 
    -- CP-element group 133: 	139 
    -- CP-element group 133: 	140 
    -- CP-element group 133: 	141 
    -- CP-element group 133: 	142 
    -- CP-element group 133: 	143 
    -- CP-element group 133: 	144 
    -- CP-element group 133: 	145 
    -- CP-element group 133: 	146 
    -- CP-element group 133: 	148 
    -- CP-element group 133: 	150 
    -- CP-element group 133: 	152 
    -- CP-element group 133:  members (112) 
      -- CP-element group 133: 	 branch_block_stmt_714/merge_stmt_1328__exit__
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460__entry__
      -- CP-element group 133: 	 branch_block_stmt_714/if_stmt_1300_if_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/if_stmt_1300_if_link/if_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/word_access_start/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/word_access_start/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/word_access_start/word_0/rr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/word_access_complete/word_0/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/word_access_start/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/word_access_start/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/word_access_start/word_0/rr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/word_access_complete/word_0/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/word_access_start/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/word_access_start/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/word_access_start/word_0/rr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/word_access_complete/word_0/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_address_resized
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_addr_resize/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_addr_resize/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_addr_resize/base_resize_req
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_addr_resize/base_resize_ack
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_plus_offset/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_plus_offset/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_plus_offset/sum_rename_req
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_base_plus_offset/sum_rename_ack
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_word_addrgen/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_word_addrgen/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_word_addrgen/root_register_req
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_word_addrgen/root_register_ack
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/word_access_start/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/word_access_start/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/word_access_start/word_0/rr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/word_access_complete/word_0/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_address_resized
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_addr_resize/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_addr_resize/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_addr_resize/base_resize_req
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_addr_resize/base_resize_ack
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_plus_offset/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_plus_offset/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_plus_offset/sum_rename_req
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_base_plus_offset/sum_rename_ack
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_word_addrgen/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_word_addrgen/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_word_addrgen/root_register_req
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_word_addrgen/root_register_ack
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/word_access_start/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/word_access_start/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/word_access_start/word_0/rr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/word_access_complete/word_0/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_update_start_
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/ifx_xelse150_whilex_xend_PhiReq/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/merge_stmt_1328_PhiReqMerge
      -- CP-element group 133: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/$entry
      -- CP-element group 133: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/$exit
      -- CP-element group 133: 	 branch_block_stmt_714/merge_stmt_1328_PhiAck/dummy
      -- 
    if_choice_transition_3934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1300_branch_ack_1, ack => zeropad3D_CP_2152_elements(133)); -- 
    rr_3959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => LOAD_col_high_1331_load_0_req_0); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => LOAD_col_high_1331_load_0_req_1); -- 
    cr_3989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1335_inst_req_1); -- 
    rr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => LOAD_pad_1344_load_0_req_0); -- 
    cr_4017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => LOAD_pad_1344_load_0_req_1); -- 
    rr_4039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => LOAD_depth_high_1347_load_0_req_0); -- 
    cr_4050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => LOAD_depth_high_1347_load_0_req_1); -- 
    rr_4089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => ptr_deref_1359_load_0_req_0); -- 
    cr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => ptr_deref_1359_load_0_req_1); -- 
    rr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => ptr_deref_1371_load_0_req_0); -- 
    cr_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => ptr_deref_1371_load_0_req_1); -- 
    cr_4169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1375_inst_req_1); -- 
    cr_4183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1379_inst_req_1); -- 
    cr_4197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(133), ack => type_cast_1418_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  place  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	841 
    -- CP-element group 134: 	842 
    -- CP-element group 134: 	844 
    -- CP-element group 134: 	845 
    -- CP-element group 134: 	846 
    -- CP-element group 134:  members (22) 
      -- CP-element group 134: 	 branch_block_stmt_714/if_stmt_1300_else_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_714/if_stmt_1300_else_link/else_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/cr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1300_branch_ack_0, ack => zeropad3D_CP_2152_elements(134)); -- 
    rr_11723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1318_inst_req_0); -- 
    cr_11728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1318_inst_req_1); -- 
    rr_11754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1310_inst_req_0); -- 
    cr_11759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(134), ack => type_cast_1310_inst_req_1); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/word_access_start/$exit
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/word_access_start/word_0/$exit
      -- CP-element group 135: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Sample/word_access_start/word_0/ra
      -- 
    ra_3960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1331_load_0_ack_0, ack => zeropad3D_CP_2152_elements(135)); -- 
    -- CP-element group 136:  fork  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	133 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136: 	149 
    -- CP-element group 136:  members (15) 
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/word_access_complete/$exit
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/word_access_complete/word_0/$exit
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/word_access_complete/word_0/ca
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/LOAD_col_high_1331_Merge/$entry
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/LOAD_col_high_1331_Merge/$exit
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/LOAD_col_high_1331_Merge/merge_req
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_col_high_1331_Update/LOAD_col_high_1331_Merge/merge_ack
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Sample/rr
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1331_load_0_ack_1, ack => zeropad3D_CP_2152_elements(136)); -- 
    rr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(136), ack => type_cast_1335_inst_req_0); -- 
    rr_4178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(136), ack => type_cast_1379_inst_req_0); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Sample/ra
      -- 
    ra_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1335_inst_ack_0, ack => zeropad3D_CP_2152_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	133 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	153 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1335_Update/ca
      -- 
    ca_3990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1335_inst_ack_1, ack => zeropad3D_CP_2152_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	133 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (5) 
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/word_access_start/$exit
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/word_access_start/word_0/$exit
      -- CP-element group 139: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Sample/word_access_start/word_0/ra
      -- 
    ra_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1344_load_0_ack_0, ack => zeropad3D_CP_2152_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	133 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	151 
    -- CP-element group 140:  members (12) 
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/word_access_complete/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/word_access_complete/word_0/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/word_access_complete/word_0/ca
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/LOAD_pad_1344_Merge/$entry
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/LOAD_pad_1344_Merge/$exit
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/LOAD_pad_1344_Merge/merge_req
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_pad_1344_Update/LOAD_pad_1344_Merge/merge_ack
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Sample/rr
      -- 
    ca_4018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1344_load_0_ack_1, ack => zeropad3D_CP_2152_elements(140)); -- 
    rr_4192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(140), ack => type_cast_1418_inst_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	133 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (5) 
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/word_access_start/$exit
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/word_access_start/word_0/$exit
      -- CP-element group 141: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Sample/word_access_start/word_0/ra
      -- 
    ra_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1347_load_0_ack_0, ack => zeropad3D_CP_2152_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	133 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	147 
    -- CP-element group 142:  members (12) 
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/word_access_complete/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/word_access_complete/word_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/word_access_complete/word_0/ca
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/LOAD_depth_high_1347_Merge/$entry
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/LOAD_depth_high_1347_Merge/$exit
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/LOAD_depth_high_1347_Merge/merge_req
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/LOAD_depth_high_1347_Update/LOAD_depth_high_1347_Merge/merge_ack
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Sample/rr
      -- 
    ca_4051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1347_load_0_ack_1, ack => zeropad3D_CP_2152_elements(142)); -- 
    rr_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(142), ack => type_cast_1375_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	133 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/word_access_start/$exit
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/word_access_start/word_0/$exit
      -- CP-element group 143: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Sample/word_access_start/word_0/ra
      -- 
    ra_4090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1359_load_0_ack_0, ack => zeropad3D_CP_2152_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	133 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	153 
    -- CP-element group 144:  members (9) 
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/word_access_complete/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/word_access_complete/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/word_access_complete/word_0/ca
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/ptr_deref_1359_Merge/$entry
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/ptr_deref_1359_Merge/$exit
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/ptr_deref_1359_Merge/merge_req
      -- CP-element group 144: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1359_Update/ptr_deref_1359_Merge/merge_ack
      -- 
    ca_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1359_load_0_ack_1, ack => zeropad3D_CP_2152_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	133 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/word_access_start/$exit
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Sample/word_access_start/word_0/ra
      -- 
    ra_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1371_load_0_ack_0, ack => zeropad3D_CP_2152_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	133 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	153 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/word_access_complete/$exit
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/ptr_deref_1371_Merge/$entry
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/ptr_deref_1371_Merge/$exit
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/ptr_deref_1371_Merge/merge_req
      -- CP-element group 146: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/ptr_deref_1371_Update/ptr_deref_1371_Merge/merge_ack
      -- 
    ca_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1371_load_0_ack_1, ack => zeropad3D_CP_2152_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	142 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Sample/ra
      -- 
    ra_4165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1375_inst_ack_0, ack => zeropad3D_CP_2152_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	133 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1375_Update/ca
      -- 
    ca_4170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1375_inst_ack_1, ack => zeropad3D_CP_2152_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	136 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Sample/ra
      -- 
    ra_4179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_0, ack => zeropad3D_CP_2152_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	133 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1379_Update/ca
      -- 
    ca_4184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_1, ack => zeropad3D_CP_2152_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	140 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Sample/ra
      -- 
    ra_4193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => zeropad3D_CP_2152_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	133 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/type_cast_1418_Update/ca
      -- 
    ca_4198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => zeropad3D_CP_2152_elements(152)); -- 
    -- CP-element group 153:  join  fork  transition  place  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	138 
    -- CP-element group 153: 	144 
    -- CP-element group 153: 	146 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	874 
    -- CP-element group 153: 	875 
    -- CP-element group 153: 	877 
    -- CP-element group 153: 	878 
    -- CP-element group 153:  members (16) 
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460__exit__
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244
      -- CP-element group 153: 	 branch_block_stmt_714/assign_stmt_1332_to_assign_stmt_1460/$exit
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Update/cr
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1469/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1476/$entry
      -- CP-element group 153: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/$entry
      -- 
    rr_11939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(153), ack => type_cast_1466_inst_req_0); -- 
    cr_11944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(153), ack => type_cast_1466_inst_req_1); -- 
    zeropad3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(138) & zeropad3D_CP_2152_elements(144) & zeropad3D_CP_2152_elements(146) & zeropad3D_CP_2152_elements(148) & zeropad3D_CP_2152_elements(150) & zeropad3D_CP_2152_elements(152);
      gj_zeropad3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	884 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Sample/ra
      -- 
    ra_4210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1487_inst_ack_0, ack => zeropad3D_CP_2152_elements(154)); -- 
    -- CP-element group 155:  branch  transition  place  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	884 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (13) 
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495__exit__
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496__entry__
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496_dead_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496_eval_test/$entry
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496_eval_test/$exit
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496_eval_test/branch_req
      -- CP-element group 155: 	 branch_block_stmt_714/R_cmp249_1497_place
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496_if_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_714/if_stmt_1496_else_link/$entry
      -- 
    ca_4215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1487_inst_ack_1, ack => zeropad3D_CP_2152_elements(155)); -- 
    branch_req_4223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(155), ack => if_stmt_1496_branch_req_0); -- 
    -- CP-element group 156:  transition  place  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	885 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_714/if_stmt_1496_if_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_714/if_stmt_1496_if_link/if_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_714/whilex_xbody244_ifx_xthen279
      -- CP-element group 156: 	 branch_block_stmt_714/whilex_xbody244_ifx_xthen279_PhiReq/$entry
      -- CP-element group 156: 	 branch_block_stmt_714/whilex_xbody244_ifx_xthen279_PhiReq/$exit
      -- 
    if_choice_transition_4228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1496_branch_ack_1, ack => zeropad3D_CP_2152_elements(156)); -- 
    -- CP-element group 157:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	161 
    -- CP-element group 157:  members (27) 
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527__entry__
      -- CP-element group 157: 	 branch_block_stmt_714/merge_stmt_1502__exit__
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1496_else_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_714/if_stmt_1496_else_link/else_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_714/whilex_xbody244_lorx_xlhsx_xfalse251
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_update_start_
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_word_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_root_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/word_access_start/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/word_access_start/word_0/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/word_access_start/word_0/rr
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/word_access_complete/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/word_access_complete/word_0/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/word_access_complete/word_0/cr
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_update_start_
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_714/whilex_xbody244_lorx_xlhsx_xfalse251_PhiReq/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/whilex_xbody244_lorx_xlhsx_xfalse251_PhiReq/$exit
      -- CP-element group 157: 	 branch_block_stmt_714/merge_stmt_1502_PhiReqMerge
      -- CP-element group 157: 	 branch_block_stmt_714/merge_stmt_1502_PhiAck/$entry
      -- CP-element group 157: 	 branch_block_stmt_714/merge_stmt_1502_PhiAck/$exit
      -- CP-element group 157: 	 branch_block_stmt_714/merge_stmt_1502_PhiAck/dummy
      -- 
    else_choice_transition_4232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1496_branch_ack_0, ack => zeropad3D_CP_2152_elements(157)); -- 
    rr_4253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(157), ack => LOAD_row_high_1504_load_0_req_0); -- 
    cr_4264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(157), ack => LOAD_row_high_1504_load_0_req_1); -- 
    cr_4283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(157), ack => type_cast_1508_inst_req_1); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (5) 
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/word_access_start/$exit
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/word_access_start/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Sample/word_access_start/word_0/ra
      -- 
    ra_4254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1504_load_0_ack_0, ack => zeropad3D_CP_2152_elements(158)); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (12) 
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/word_access_complete/$exit
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/word_access_complete/word_0/$exit
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/word_access_complete/word_0/ca
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/LOAD_row_high_1504_Merge/$entry
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/LOAD_row_high_1504_Merge/$exit
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/LOAD_row_high_1504_Merge/merge_req
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/LOAD_row_high_1504_Update/LOAD_row_high_1504_Merge/merge_ack
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Sample/rr
      -- 
    ca_4265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1504_load_0_ack_1, ack => zeropad3D_CP_2152_elements(159)); -- 
    rr_4278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(159), ack => type_cast_1508_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Sample/ra
      -- 
    ra_4279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1508_inst_ack_0, ack => zeropad3D_CP_2152_elements(160)); -- 
    -- CP-element group 161:  branch  transition  place  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	157 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (13) 
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528__entry__
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527__exit__
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/$exit
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_714/assign_stmt_1505_to_assign_stmt_1527/type_cast_1508_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528_dead_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528_eval_test/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528_eval_test/$exit
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528_eval_test/branch_req
      -- CP-element group 161: 	 branch_block_stmt_714/R_cmp260_1529_place
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528_if_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_714/if_stmt_1528_else_link/$entry
      -- 
    ca_4284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1508_inst_ack_1, ack => zeropad3D_CP_2152_elements(161)); -- 
    branch_req_4292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(161), ack => if_stmt_1528_branch_req_0); -- 
    -- CP-element group 162:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: 	165 
    -- CP-element group 162:  members (18) 
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546__entry__
      -- CP-element group 162: 	 branch_block_stmt_714/merge_stmt_1534__exit__
      -- CP-element group 162: 	 branch_block_stmt_714/if_stmt_1528_if_link/$exit
      -- CP-element group 162: 	 branch_block_stmt_714/if_stmt_1528_if_link/if_choice_transition
      -- CP-element group 162: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_lorx_xlhsx_xfalse262
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/$entry
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_update_start_
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Update/cr
      -- CP-element group 162: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_lorx_xlhsx_xfalse262_PhiReq/$entry
      -- CP-element group 162: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_lorx_xlhsx_xfalse262_PhiReq/$exit
      -- CP-element group 162: 	 branch_block_stmt_714/merge_stmt_1534_PhiReqMerge
      -- CP-element group 162: 	 branch_block_stmt_714/merge_stmt_1534_PhiAck/$entry
      -- CP-element group 162: 	 branch_block_stmt_714/merge_stmt_1534_PhiAck/$exit
      -- CP-element group 162: 	 branch_block_stmt_714/merge_stmt_1534_PhiAck/dummy
      -- 
    if_choice_transition_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1528_branch_ack_1, ack => zeropad3D_CP_2152_elements(162)); -- 
    rr_4314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(162), ack => type_cast_1538_inst_req_0); -- 
    cr_4319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(162), ack => type_cast_1538_inst_req_1); -- 
    -- CP-element group 163:  transition  place  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	885 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_714/if_stmt_1528_else_link/$exit
      -- CP-element group 163: 	 branch_block_stmt_714/if_stmt_1528_else_link/else_choice_transition
      -- CP-element group 163: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_ifx_xthen279
      -- CP-element group 163: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_ifx_xthen279_PhiReq/$entry
      -- CP-element group 163: 	 branch_block_stmt_714/lorx_xlhsx_xfalse251_ifx_xthen279_PhiReq/$exit
      -- 
    else_choice_transition_4301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1528_branch_ack_0, ack => zeropad3D_CP_2152_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Sample/ra
      -- 
    ra_4315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_0, ack => zeropad3D_CP_2152_elements(164)); -- 
    -- CP-element group 165:  branch  transition  place  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546__exit__
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547__entry__
      -- CP-element group 165: 	 branch_block_stmt_714/R_cmp267_1548_place
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547_else_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547_if_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/assign_stmt_1539_to_assign_stmt_1546/type_cast_1538_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547_dead_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547_eval_test/$entry
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547_eval_test/$exit
      -- CP-element group 165: 	 branch_block_stmt_714/if_stmt_1547_eval_test/branch_req
      -- 
    ca_4320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_1, ack => zeropad3D_CP_2152_elements(165)); -- 
    branch_req_4328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(165), ack => if_stmt_1547_branch_req_0); -- 
    -- CP-element group 166:  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	885 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_ifx_xthen279
      -- CP-element group 166: 	 branch_block_stmt_714/if_stmt_1547_if_link/if_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_714/if_stmt_1547_if_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_ifx_xthen279_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_ifx_xthen279_PhiReq/$exit
      -- 
    if_choice_transition_4333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1547_branch_ack_1, ack => zeropad3D_CP_2152_elements(166)); -- 
    -- CP-element group 167:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: 	169 
    -- CP-element group 167: 	171 
    -- CP-element group 167:  members (27) 
      -- CP-element group 167: 	 branch_block_stmt_714/merge_stmt_1553__exit__
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572__entry__
      -- CP-element group 167: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_lorx_xlhsx_xfalse269
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_update_start_
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/word_access_complete/word_0/cr
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/word_access_complete/word_0/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/word_access_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/word_access_start/word_0/rr
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/word_access_start/word_0/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1547_else_link/else_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/word_access_start/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_root_address_calculated
      -- CP-element group 167: 	 branch_block_stmt_714/if_stmt_1547_else_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_word_address_calculated
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_update_start_
      -- CP-element group 167: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_lorx_xlhsx_xfalse269_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/lorx_xlhsx_xfalse262_lorx_xlhsx_xfalse269_PhiReq/$exit
      -- CP-element group 167: 	 branch_block_stmt_714/merge_stmt_1553_PhiReqMerge
      -- CP-element group 167: 	 branch_block_stmt_714/merge_stmt_1553_PhiAck/$entry
      -- CP-element group 167: 	 branch_block_stmt_714/merge_stmt_1553_PhiAck/$exit
      -- CP-element group 167: 	 branch_block_stmt_714/merge_stmt_1553_PhiAck/dummy
      -- 
    else_choice_transition_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1547_branch_ack_0, ack => zeropad3D_CP_2152_elements(167)); -- 
    cr_4369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(167), ack => LOAD_col_high_1555_load_0_req_1); -- 
    rr_4358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(167), ack => LOAD_col_high_1555_load_0_req_0); -- 
    cr_4388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(167), ack => type_cast_1559_inst_req_1); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (5) 
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/word_access_start/word_0/ra
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/word_access_start/word_0/$exit
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/word_access_start/$exit
      -- CP-element group 168: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Sample/$exit
      -- 
    ra_4359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1555_load_0_ack_0, ack => zeropad3D_CP_2152_elements(168)); -- 
    -- CP-element group 169:  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (12) 
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/LOAD_col_high_1555_Merge/merge_ack
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/LOAD_col_high_1555_Merge/merge_req
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/LOAD_col_high_1555_Merge/$exit
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/LOAD_col_high_1555_Merge/$entry
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/word_access_complete/word_0/ca
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/word_access_complete/word_0/$exit
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/word_access_complete/$exit
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/LOAD_col_high_1555_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Sample/rr
      -- CP-element group 169: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Sample/$entry
      -- 
    ca_4370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1555_load_0_ack_1, ack => zeropad3D_CP_2152_elements(169)); -- 
    rr_4383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(169), ack => type_cast_1559_inst_req_0); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_sample_completed_
      -- 
    ra_4384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_0, ack => zeropad3D_CP_2152_elements(170)); -- 
    -- CP-element group 171:  branch  transition  place  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	167 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (13) 
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572__exit__
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573__entry__
      -- CP-element group 171: 	 branch_block_stmt_714/R_cmp277_1574_place
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/$exit
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573_else_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573_if_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573_eval_test/branch_req
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573_eval_test/$exit
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573_eval_test/$entry
      -- CP-element group 171: 	 branch_block_stmt_714/if_stmt_1573_dead_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_714/assign_stmt_1556_to_assign_stmt_1572/type_cast_1559_update_completed_
      -- 
    ca_4389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_1, ack => zeropad3D_CP_2152_elements(171)); -- 
    branch_req_4397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(171), ack => if_stmt_1573_branch_req_0); -- 
    -- CP-element group 172:  fork  transition  place  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	188 
    -- CP-element group 172: 	189 
    -- CP-element group 172: 	191 
    -- CP-element group 172: 	193 
    -- CP-element group 172: 	195 
    -- CP-element group 172: 	197 
    -- CP-element group 172: 	199 
    -- CP-element group 172: 	201 
    -- CP-element group 172: 	203 
    -- CP-element group 172: 	206 
    -- CP-element group 172:  members (46) 
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742__entry__
      -- CP-element group 172: 	 branch_block_stmt_714/merge_stmt_1637__exit__
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_complete/req
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_update_start
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_update_start
      -- CP-element group 172: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xelse300
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Update/req
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/if_stmt_1573_if_link/if_choice_transition
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Update/req
      -- CP-element group 172: 	 branch_block_stmt_714/if_stmt_1573_if_link/$exit
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_update_start_
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_complete/req
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xelse300_PhiReq/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xelse300_PhiReq/$exit
      -- CP-element group 172: 	 branch_block_stmt_714/merge_stmt_1637_PhiReqMerge
      -- CP-element group 172: 	 branch_block_stmt_714/merge_stmt_1637_PhiAck/$entry
      -- CP-element group 172: 	 branch_block_stmt_714/merge_stmt_1637_PhiAck/$exit
      -- CP-element group 172: 	 branch_block_stmt_714/merge_stmt_1637_PhiAck/dummy
      -- 
    if_choice_transition_4402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1573_branch_ack_1, ack => zeropad3D_CP_2152_elements(172)); -- 
    rr_4560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => type_cast_1641_inst_req_0); -- 
    req_4735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => addr_of_1737_final_reg_req_1); -- 
    cr_4689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => type_cast_1730_inst_req_1); -- 
    req_4720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => array_obj_ref_1736_index_offset_req_1); -- 
    cr_4670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => ptr_deref_1716_load_0_req_1); -- 
    req_4610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => array_obj_ref_1711_index_offset_req_1); -- 
    cr_4579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => type_cast_1705_inst_req_1); -- 
    cr_4565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => type_cast_1641_inst_req_1); -- 
    req_4625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => addr_of_1712_final_reg_req_1); -- 
    cr_4785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(172), ack => ptr_deref_1740_store_0_req_1); -- 
    -- CP-element group 173:  transition  place  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	885 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xthen279
      -- CP-element group 173: 	 branch_block_stmt_714/if_stmt_1573_else_link/else_choice_transition
      -- CP-element group 173: 	 branch_block_stmt_714/if_stmt_1573_else_link/$exit
      -- CP-element group 173: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xthen279_PhiReq/$entry
      -- CP-element group 173: 	 branch_block_stmt_714/lorx_xlhsx_xfalse269_ifx_xthen279_PhiReq/$exit
      -- 
    else_choice_transition_4406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1573_branch_ack_0, ack => zeropad3D_CP_2152_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	885 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Sample/$exit
      -- 
    ra_4420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_0, ack => zeropad3D_CP_2152_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	885 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Update/$exit
      -- 
    ca_4425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_1, ack => zeropad3D_CP_2152_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	885 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Sample/ra
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_sample_completed_
      -- 
    ra_4434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1588_inst_ack_0, ack => zeropad3D_CP_2152_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	885 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Update/ca
      -- CP-element group 177: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_update_completed_
      -- 
    ca_4439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1588_inst_ack_1, ack => zeropad3D_CP_2152_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_sample_start_
      -- 
    rr_4447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(178), ack => type_cast_1622_inst_req_0); -- 
    zeropad3D_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(175) & zeropad3D_CP_2152_elements(177);
      gj_zeropad3D_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_sample_completed_
      -- 
    ra_4448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1622_inst_ack_0, ack => zeropad3D_CP_2152_elements(179)); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	885 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (16) 
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Sample/req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_scale_1/scale_rename_ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_scale_1/scale_rename_req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_scale_1/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_scale_1/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_resize_1/index_resize_ack
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_resize_1/index_resize_req
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_resize_1/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_resize_1/$entry
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_computed_1
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_scaled_1
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_index_resized_1
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_update_completed_
      -- 
    ca_4453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1622_inst_ack_1, ack => zeropad3D_CP_2152_elements(180)); -- 
    req_4478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(180), ack => array_obj_ref_1628_index_offset_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	187 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Sample/ack
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_sample_complete
      -- 
    ack_4479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1628_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	885 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (11) 
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Update/ack
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_offset_calculated
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_root_address_calculated
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_request/req
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_request/$entry
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_base_plus_offset/sum_rename_ack
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_base_plus_offset/sum_rename_req
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_base_plus_offset/$exit
      -- CP-element group 182: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_base_plus_offset/$entry
      -- 
    ack_4484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1628_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(182)); -- 
    req_4493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(182), ack => addr_of_1629_final_reg_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_request/ack
      -- CP-element group 183: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_request/$exit
      -- 
    ack_4494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1629_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(183)); -- 
    -- CP-element group 184:  join  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	885 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (28) 
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_addr_resize/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_addr_resize/$exit
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_address_resized
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_root_address_calculated
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_word_address_calculated
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_address_calculated
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_complete/ack
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/word_access_start/word_0/rr
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/word_access_start/word_0/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_complete/$exit
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/word_access_start/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/ptr_deref_1632_Split/split_ack
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/ptr_deref_1632_Split/split_req
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/ptr_deref_1632_Split/$exit
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/ptr_deref_1632_Split/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_word_addrgen/root_register_ack
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_word_addrgen/root_register_req
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_word_addrgen/$exit
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_word_addrgen/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_plus_offset/sum_rename_ack
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_plus_offset/sum_rename_req
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_plus_offset/$exit
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_plus_offset/$entry
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_addr_resize/base_resize_ack
      -- CP-element group 184: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_base_addr_resize/base_resize_req
      -- 
    ack_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1629_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(184)); -- 
    rr_4537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(184), ack => ptr_deref_1632_store_0_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (5) 
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/word_access_start/word_0/ra
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/word_access_start/word_0/$exit
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/word_access_start/$exit
      -- CP-element group 185: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Sample/$exit
      -- 
    ra_4538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1632_store_0_ack_0, ack => zeropad3D_CP_2152_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	885 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (5) 
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/word_access_complete/word_0/ca
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/word_access_complete/word_0/$exit
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/word_access_complete/$exit
      -- CP-element group 186: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/$exit
      -- 
    ca_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1632_store_0_ack_1, ack => zeropad3D_CP_2152_elements(186)); -- 
    -- CP-element group 187:  join  transition  place  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	181 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	886 
    -- CP-element group 187:  members (5) 
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635__exit__
      -- CP-element group 187: 	 branch_block_stmt_714/ifx_xthen279_ifx_xend348
      -- CP-element group 187: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/$exit
      -- CP-element group 187: 	 branch_block_stmt_714/ifx_xthen279_ifx_xend348_PhiReq/$entry
      -- CP-element group 187: 	 branch_block_stmt_714/ifx_xthen279_ifx_xend348_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(181) & zeropad3D_CP_2152_elements(186);
      gj_zeropad3D_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	172 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Sample/ra
      -- CP-element group 188: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_sample_completed_
      -- 
    ra_4561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1641_inst_ack_0, ack => zeropad3D_CP_2152_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	172 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189: 	198 
    -- CP-element group 189:  members (9) 
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1641_Update/$exit
      -- 
    ca_4566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1641_inst_ack_1, ack => zeropad3D_CP_2152_elements(189)); -- 
    rr_4574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(189), ack => type_cast_1705_inst_req_0); -- 
    rr_4684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(189), ack => type_cast_1730_inst_req_0); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_sample_completed_
      -- 
    ra_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1705_inst_ack_0, ack => zeropad3D_CP_2152_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	172 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (16) 
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Sample/req
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_scale_1/scale_rename_ack
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_scale_1/scale_rename_req
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_scale_1/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_scale_1/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_resize_1/index_resize_ack
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_resize_1/index_resize_req
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_resize_1/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_resize_1/$entry
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_computed_1
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_scaled_1
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_index_resized_1
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1705_update_completed_
      -- 
    ca_4580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1705_inst_ack_1, ack => zeropad3D_CP_2152_elements(191)); -- 
    req_4605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(191), ack => array_obj_ref_1711_index_offset_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	207 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Sample/ack
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_sample_complete
      -- 
    ack_4606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1711_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	172 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (11) 
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_base_plus_offset/sum_rename_ack
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_request/req
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_base_plus_offset/sum_rename_req
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_base_plus_offset/$exit
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_base_plus_offset/$entry
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Update/ack
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_offset_calculated
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_root_address_calculated
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_request/$entry
      -- CP-element group 193: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1711_final_index_sum_regn_Update/$exit
      -- 
    ack_4611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1711_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(193)); -- 
    req_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(193), ack => addr_of_1712_final_reg_req_0); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_request/ack
      -- CP-element group 194: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_request/$exit
      -- CP-element group 194: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_sample_completed_
      -- 
    ack_4621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1712_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(194)); -- 
    -- CP-element group 195:  join  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	172 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (24) 
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_complete/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/word_access_start/word_0/rr
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/word_access_start/word_0/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/word_access_start/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_word_addrgen/root_register_ack
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_word_addrgen/root_register_req
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_word_addrgen/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_word_addrgen/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_plus_offset/sum_rename_ack
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_plus_offset/sum_rename_req
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_plus_offset/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_plus_offset/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_addr_resize/base_resize_ack
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_addr_resize/base_resize_req
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_addr_resize/$exit
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_addr_resize/$entry
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_address_resized
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_root_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_word_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_base_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1712_complete/ack
      -- 
    ack_4626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1712_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(195)); -- 
    rr_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(195), ack => ptr_deref_1716_load_0_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (5) 
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/word_access_start/word_0/ra
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/word_access_start/word_0/$exit
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/word_access_start/$exit
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_sample_completed_
      -- 
    ra_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1716_load_0_ack_0, ack => zeropad3D_CP_2152_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	172 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	204 
    -- CP-element group 197:  members (9) 
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/ptr_deref_1716_Merge/merge_ack
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/ptr_deref_1716_Merge/merge_req
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/ptr_deref_1716_Merge/$exit
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/ptr_deref_1716_Merge/$entry
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/word_access_complete/word_0/ca
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/word_access_complete/word_0/$exit
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1716_Update/word_access_complete/$exit
      -- 
    ca_4671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1716_load_0_ack_1, ack => zeropad3D_CP_2152_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	189 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Sample/$exit
      -- 
    ra_4685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1730_inst_ack_0, ack => zeropad3D_CP_2152_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	172 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (16) 
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_resize_1/index_resize_ack
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_scale_1/$entry
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_resize_1/index_resize_req
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_scale_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_resize_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_resize_1/$entry
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_computed_1
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_scaled_1
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_resized_1
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Sample/req
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_scale_1/scale_rename_ack
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/type_cast_1730_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_index_scale_1/scale_rename_req
      -- 
    ca_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1730_inst_ack_1, ack => zeropad3D_CP_2152_elements(199)); -- 
    req_4715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(199), ack => array_obj_ref_1736_index_offset_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	207 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Sample/ack
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_sample_complete
      -- 
    ack_4716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	172 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (11) 
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_base_plus_offset/$exit
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_base_plus_offset/$entry
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_offset_calculated
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_root_address_calculated
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_request/req
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Update/ack
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_base_plus_offset/sum_rename_ack
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_base_plus_offset/sum_rename_req
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_request/$entry
      -- CP-element group 201: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/array_obj_ref_1736_final_index_sum_regn_Update/$exit
      -- 
    ack_4721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(201)); -- 
    req_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(201), ack => addr_of_1737_final_reg_req_0); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_request/ack
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_request/$exit
      -- 
    ack_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1737_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	172 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (19) 
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_word_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_root_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_complete/$exit
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/addr_of_1737_complete/ack
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_address_resized
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_addr_resize/$entry
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_addr_resize/$exit
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_addr_resize/base_resize_req
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_addr_resize/base_resize_ack
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_plus_offset/$entry
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_plus_offset/$exit
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_plus_offset/sum_rename_req
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_base_plus_offset/sum_rename_ack
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_word_addrgen/$entry
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_word_addrgen/$exit
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_word_addrgen/root_register_req
      -- CP-element group 203: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_word_addrgen/root_register_ack
      -- 
    ack_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1737_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	197 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (9) 
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/ptr_deref_1740_Split/$entry
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/ptr_deref_1740_Split/$exit
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/ptr_deref_1740_Split/split_req
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/ptr_deref_1740_Split/split_ack
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/word_access_start/$entry
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/word_access_start/word_0/$entry
      -- CP-element group 204: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/word_access_start/word_0/rr
      -- 
    rr_4774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(204), ack => ptr_deref_1740_store_0_req_0); -- 
    zeropad3D_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(197) & zeropad3D_CP_2152_elements(203);
      gj_zeropad3D_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/word_access_start/$exit
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/word_access_start/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Sample/word_access_start/word_0/ra
      -- 
    ra_4775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1740_store_0_ack_0, ack => zeropad3D_CP_2152_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	172 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/word_access_complete/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/word_access_complete/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/ptr_deref_1740_Update/word_access_complete/word_0/ca
      -- 
    ca_4786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1740_store_0_ack_1, ack => zeropad3D_CP_2152_elements(206)); -- 
    -- CP-element group 207:  join  transition  place  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	192 
    -- CP-element group 207: 	200 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	886 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742__exit__
      -- CP-element group 207: 	 branch_block_stmt_714/ifx_xelse300_ifx_xend348
      -- CP-element group 207: 	 branch_block_stmt_714/assign_stmt_1642_to_assign_stmt_1742/$exit
      -- CP-element group 207: 	 branch_block_stmt_714/ifx_xelse300_ifx_xend348_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_714/ifx_xelse300_ifx_xend348_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(192) & zeropad3D_CP_2152_elements(200) & zeropad3D_CP_2152_elements(206);
      gj_zeropad3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	886 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Sample/ra
      -- 
    ra_4798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_0, ack => zeropad3D_CP_2152_elements(208)); -- 
    -- CP-element group 209:  branch  transition  place  input  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	886 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762__exit__
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763__entry__
      -- CP-element group 209: 	 branch_block_stmt_714/R_cmp356_1764_place
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/$exit
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Update/ca
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763_eval_test/branch_req
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_714/if_stmt_1763_else_link/$entry
      -- 
    ca_4803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_1, ack => zeropad3D_CP_2152_elements(209)); -- 
    branch_req_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(209), ack => if_stmt_1763_branch_req_0); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	895 
    -- CP-element group 210: 	896 
    -- CP-element group 210: 	898 
    -- CP-element group 210: 	899 
    -- CP-element group 210: 	901 
    -- CP-element group 210: 	902 
    -- CP-element group 210:  members (40) 
      -- CP-element group 210: 	 branch_block_stmt_714/merge_stmt_1769__exit__
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1775__entry__
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1775__exit__
      -- CP-element group 210: 	 branch_block_stmt_714/if_stmt_1763_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/if_stmt_1763_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xend348_ifx_xthen358
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1775/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/assign_stmt_1775/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xend348_ifx_xthen358_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xend348_ifx_xthen358_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/merge_stmt_1769_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_714/merge_stmt_1769_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/merge_stmt_1769_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_714/merge_stmt_1769_PhiAck/dummy
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1763_branch_ack_1, ack => zeropad3D_CP_2152_elements(210)); -- 
    rr_12145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(210), ack => type_cast_1871_inst_req_0); -- 
    cr_12150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(210), ack => type_cast_1871_inst_req_1); -- 
    rr_12168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(210), ack => type_cast_1865_inst_req_0); -- 
    cr_12173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(210), ack => type_cast_1865_inst_req_1); -- 
    rr_12191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(210), ack => type_cast_1859_inst_req_0); -- 
    cr_12196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(210), ack => type_cast_1859_inst_req_1); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211: 	213 
    -- CP-element group 211: 	214 
    -- CP-element group 211: 	215 
    -- CP-element group 211: 	217 
    -- CP-element group 211: 	220 
    -- CP-element group 211: 	222 
    -- CP-element group 211: 	223 
    -- CP-element group 211: 	224 
    -- CP-element group 211: 	226 
    -- CP-element group 211:  members (54) 
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848__entry__
      -- CP-element group 211: 	 branch_block_stmt_714/merge_stmt_1777__exit__
      -- CP-element group 211: 	 branch_block_stmt_714/if_stmt_1763_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/if_stmt_1763_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_714/ifx_xend348_ifx_xelse363
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_word_address_calculated
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_root_address_calculated
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/word_access_start/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/word_access_start/word_0/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/word_access_start/word_0/rr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/word_access_complete/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/word_access_complete/word_0/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/word_access_complete/word_0/cr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_word_address_calculated
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_root_address_calculated
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/word_access_start/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/word_access_start/word_0/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/word_access_start/word_0/rr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/word_access_complete/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/word_access_complete/word_0/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/word_access_complete/word_0/cr
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_update_start_
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_714/ifx_xend348_ifx_xelse363_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/ifx_xend348_ifx_xelse363_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/merge_stmt_1777_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_714/merge_stmt_1777_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_714/merge_stmt_1777_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_714/merge_stmt_1777_PhiAck/dummy
      -- 
    else_choice_transition_4820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1763_branch_ack_0, ack => zeropad3D_CP_2152_elements(211)); -- 
    rr_4836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1787_inst_req_0); -- 
    cr_4841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1787_inst_req_1); -- 
    rr_4858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => LOAD_col_high_1790_load_0_req_0); -- 
    cr_4869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => LOAD_col_high_1790_load_0_req_1); -- 
    cr_4888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1794_inst_req_1); -- 
    cr_4902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1808_inst_req_1); -- 
    cr_4916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1824_inst_req_1); -- 
    rr_4933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => LOAD_row_high_1827_load_0_req_0); -- 
    cr_4944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => LOAD_row_high_1827_load_0_req_1); -- 
    cr_4963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(211), ack => type_cast_1831_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Sample/ra
      -- 
    ra_4837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1787_inst_ack_0, ack => zeropad3D_CP_2152_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	218 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1787_Update/ca
      -- 
    ca_4842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1787_inst_ack_1, ack => zeropad3D_CP_2152_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	211 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (5) 
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/word_access_start/$exit
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/word_access_start/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Sample/word_access_start/word_0/ra
      -- 
    ra_4859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1790_load_0_ack_0, ack => zeropad3D_CP_2152_elements(214)); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	211 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (12) 
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/word_access_complete/$exit
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/word_access_complete/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/word_access_complete/word_0/ca
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/LOAD_col_high_1790_Merge/$entry
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/LOAD_col_high_1790_Merge/$exit
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/LOAD_col_high_1790_Merge/merge_req
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_col_high_1790_Update/LOAD_col_high_1790_Merge/merge_ack
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Sample/rr
      -- 
    ca_4870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1790_load_0_ack_1, ack => zeropad3D_CP_2152_elements(215)); -- 
    rr_4883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(215), ack => type_cast_1794_inst_req_0); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Sample/ra
      -- 
    ra_4884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1794_inst_ack_0, ack => zeropad3D_CP_2152_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	211 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1794_Update/ca
      -- 
    ca_4889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1794_inst_ack_1, ack => zeropad3D_CP_2152_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	213 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Sample/rr
      -- 
    rr_4897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(218), ack => type_cast_1808_inst_req_0); -- 
    zeropad3D_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(213) & zeropad3D_CP_2152_elements(217);
      gj_zeropad3D_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Sample/ra
      -- 
    ra_4898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_0, ack => zeropad3D_CP_2152_elements(219)); -- 
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	211 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1808_Update/ca
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Sample/rr
      -- 
    ca_4903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_1, ack => zeropad3D_CP_2152_elements(220)); -- 
    rr_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(220), ack => type_cast_1824_inst_req_0); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Sample/ra
      -- 
    ra_4912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1824_inst_ack_0, ack => zeropad3D_CP_2152_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	211 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	227 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1824_Update/ca
      -- 
    ca_4917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1824_inst_ack_1, ack => zeropad3D_CP_2152_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	211 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (5) 
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/word_access_start/$exit
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/word_access_start/word_0/$exit
      -- CP-element group 223: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Sample/word_access_start/word_0/ra
      -- 
    ra_4934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1827_load_0_ack_0, ack => zeropad3D_CP_2152_elements(223)); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	211 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (12) 
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/word_access_complete/$exit
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/word_access_complete/word_0/$exit
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/word_access_complete/word_0/ca
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/LOAD_row_high_1827_Merge/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/LOAD_row_high_1827_Merge/$exit
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/LOAD_row_high_1827_Merge/merge_req
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/LOAD_row_high_1827_Update/LOAD_row_high_1827_Merge/merge_ack
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_sample_start_
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Sample/rr
      -- 
    ca_4945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1827_load_0_ack_1, ack => zeropad3D_CP_2152_elements(224)); -- 
    rr_4958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(224), ack => type_cast_1831_inst_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Sample/ra
      -- 
    ra_4959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_0, ack => zeropad3D_CP_2152_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	211 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/type_cast_1831_Update/ca
      -- 
    ca_4964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_1, ack => zeropad3D_CP_2152_elements(226)); -- 
    -- CP-element group 227:  branch  join  transition  place  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	222 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (10) 
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849__entry__
      -- CP-element group 227: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848__exit__
      -- CP-element group 227: 	 branch_block_stmt_714/assign_stmt_1783_to_assign_stmt_1848/$exit
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849_dead_link/$entry
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849_eval_test/$entry
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849_eval_test/$exit
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849_eval_test/branch_req
      -- CP-element group 227: 	 branch_block_stmt_714/R_cmp390_1850_place
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849_if_link/$entry
      -- CP-element group 227: 	 branch_block_stmt_714/if_stmt_1849_else_link/$entry
      -- 
    branch_req_4972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(227), ack => if_stmt_1849_branch_req_0); -- 
    zeropad3D_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(222) & zeropad3D_CP_2152_elements(226);
      gj_zeropad3D_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: 	231 
    -- CP-element group 228: 	233 
    -- CP-element group 228: 	234 
    -- CP-element group 228: 	235 
    -- CP-element group 228: 	236 
    -- CP-element group 228: 	237 
    -- CP-element group 228: 	238 
    -- CP-element group 228: 	239 
    -- CP-element group 228: 	240 
    -- CP-element group 228: 	241 
    -- CP-element group 228: 	242 
    -- CP-element group 228: 	243 
    -- CP-element group 228: 	245 
    -- CP-element group 228: 	247 
    -- CP-element group 228: 	249 
    -- CP-element group 228:  members (124) 
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012__entry__
      -- CP-element group 228: 	 branch_block_stmt_714/merge_stmt_1877__exit__
      -- CP-element group 228: 	 branch_block_stmt_714/if_stmt_1849_if_link/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/if_stmt_1849_if_link/if_choice_transition
      -- CP-element group 228: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_word_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_root_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/word_access_start/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/word_access_start/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/word_access_start/word_0/rr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_word_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_root_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/word_access_start/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/word_access_start/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/word_access_start/word_0/rr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_word_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_root_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/word_access_start/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/word_access_start/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/word_access_start/word_0/rr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_word_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_root_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/word_access_start/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/word_access_start/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/word_access_start/word_0/rr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_word_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_root_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_address_resized
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_addr_resize/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_addr_resize/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_addr_resize/base_resize_req
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_addr_resize/base_resize_ack
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_plus_offset/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_plus_offset/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_plus_offset/sum_rename_req
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_base_plus_offset/sum_rename_ack
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_word_addrgen/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_word_addrgen/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_word_addrgen/root_register_req
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_word_addrgen/root_register_ack
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/word_access_start/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/word_access_start/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/word_access_start/word_0/rr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_word_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_root_address_calculated
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_address_resized
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_addr_resize/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_addr_resize/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_addr_resize/base_resize_req
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_addr_resize/base_resize_ack
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_plus_offset/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_plus_offset/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_plus_offset/sum_rename_req
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_base_plus_offset/sum_rename_ack
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_word_addrgen/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_word_addrgen/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_word_addrgen/root_register_req
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_word_addrgen/root_register_ack
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/word_access_start/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/word_access_start/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/word_access_start/word_0/rr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/word_access_complete/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/word_access_complete/word_0/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/word_access_complete/word_0/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_update_start_
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/ifx_xelse363_whilex_xend400_PhiReq/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/merge_stmt_1877_PhiReqMerge
      -- CP-element group 228: 	 branch_block_stmt_714/merge_stmt_1877_PhiAck/$entry
      -- CP-element group 228: 	 branch_block_stmt_714/merge_stmt_1877_PhiAck/$exit
      -- CP-element group 228: 	 branch_block_stmt_714/merge_stmt_1877_PhiAck/dummy
      -- 
    if_choice_transition_4977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1849_branch_ack_1, ack => zeropad3D_CP_2152_elements(228)); -- 
    rr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_row_high_1880_load_0_req_0); -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_row_high_1880_load_0_req_1); -- 
    cr_5032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => type_cast_1884_inst_req_1); -- 
    rr_5049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_pad_1893_load_0_req_0); -- 
    cr_5060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_pad_1893_load_0_req_1); -- 
    rr_5082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_depth_high_1896_load_0_req_0); -- 
    cr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_depth_high_1896_load_0_req_1); -- 
    rr_5115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_col_high_1899_load_0_req_0); -- 
    cr_5126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => LOAD_col_high_1899_load_0_req_1); -- 
    rr_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => ptr_deref_1911_load_0_req_0); -- 
    cr_5176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => ptr_deref_1911_load_0_req_1); -- 
    rr_5215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => ptr_deref_1923_load_0_req_0); -- 
    cr_5226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => ptr_deref_1923_load_0_req_1); -- 
    cr_5245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => type_cast_1927_inst_req_1); -- 
    cr_5259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => type_cast_1931_inst_req_1); -- 
    cr_5273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(228), ack => type_cast_1970_inst_req_1); -- 
    -- CP-element group 229:  fork  transition  place  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	887 
    -- CP-element group 229: 	888 
    -- CP-element group 229: 	889 
    -- CP-element group 229: 	891 
    -- CP-element group 229: 	892 
    -- CP-element group 229:  members (22) 
      -- CP-element group 229: 	 branch_block_stmt_714/if_stmt_1849_else_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_714/if_stmt_1849_else_link/else_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1868/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Update/cr
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1849_branch_ack_0, ack => zeropad3D_CP_2152_elements(229)); -- 
    rr_12096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(229), ack => type_cast_1867_inst_req_0); -- 
    cr_12101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(229), ack => type_cast_1867_inst_req_1); -- 
    rr_12119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(229), ack => type_cast_1861_inst_req_0); -- 
    cr_12124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(229), ack => type_cast_1861_inst_req_1); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Sample/word_access_start/word_0/ra
      -- 
    ra_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1880_load_0_ack_0, ack => zeropad3D_CP_2152_elements(230)); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	228 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (12) 
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/word_access_complete/word_0/ca
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/LOAD_row_high_1880_Merge/$entry
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/LOAD_row_high_1880_Merge/$exit
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/LOAD_row_high_1880_Merge/merge_req
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_row_high_1880_Update/LOAD_row_high_1880_Merge/merge_ack
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Sample/rr
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_1880_load_0_ack_1, ack => zeropad3D_CP_2152_elements(231)); -- 
    rr_5027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(231), ack => type_cast_1884_inst_req_0); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Sample/ra
      -- 
    ra_5028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1884_inst_ack_0, ack => zeropad3D_CP_2152_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	228 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	250 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1884_Update/ca
      -- 
    ca_5033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1884_inst_ack_1, ack => zeropad3D_CP_2152_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	228 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (5) 
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/word_access_start/$exit
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/word_access_start/word_0/$exit
      -- CP-element group 234: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Sample/word_access_start/word_0/ra
      -- 
    ra_5050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1893_load_0_ack_0, ack => zeropad3D_CP_2152_elements(234)); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	228 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	248 
    -- CP-element group 235:  members (12) 
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/word_access_complete/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/word_access_complete/word_0/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/word_access_complete/word_0/ca
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/LOAD_pad_1893_Merge/$entry
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/LOAD_pad_1893_Merge/$exit
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/LOAD_pad_1893_Merge/merge_req
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_pad_1893_Update/LOAD_pad_1893_Merge/merge_ack
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Sample/rr
      -- 
    ca_5061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1893_load_0_ack_1, ack => zeropad3D_CP_2152_elements(235)); -- 
    rr_5268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(235), ack => type_cast_1970_inst_req_0); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	228 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/word_access_start/$exit
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/word_access_start/word_0/$exit
      -- CP-element group 236: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Sample/word_access_start/word_0/ra
      -- 
    ra_5083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1896_load_0_ack_0, ack => zeropad3D_CP_2152_elements(236)); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	228 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	244 
    -- CP-element group 237:  members (12) 
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/word_access_complete/$exit
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/word_access_complete/word_0/$exit
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/word_access_complete/word_0/ca
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/LOAD_depth_high_1896_Merge/$entry
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/LOAD_depth_high_1896_Merge/$exit
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/LOAD_depth_high_1896_Merge/merge_req
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_depth_high_1896_Update/LOAD_depth_high_1896_Merge/merge_ack
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Sample/rr
      -- 
    ca_5094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_1896_load_0_ack_1, ack => zeropad3D_CP_2152_elements(237)); -- 
    rr_5240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(237), ack => type_cast_1927_inst_req_0); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	228 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (5) 
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/word_access_start/$exit
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/word_access_start/word_0/$exit
      -- CP-element group 238: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Sample/word_access_start/word_0/ra
      -- 
    ra_5116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1899_load_0_ack_0, ack => zeropad3D_CP_2152_elements(238)); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	228 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	246 
    -- CP-element group 239:  members (12) 
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/word_access_complete/$exit
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/word_access_complete/word_0/$exit
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/word_access_complete/word_0/ca
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/LOAD_col_high_1899_Merge/$entry
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/LOAD_col_high_1899_Merge/$exit
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/LOAD_col_high_1899_Merge/merge_req
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/LOAD_col_high_1899_Update/LOAD_col_high_1899_Merge/merge_ack
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Sample/rr
      -- 
    ca_5127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_1899_load_0_ack_1, ack => zeropad3D_CP_2152_elements(239)); -- 
    rr_5254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(239), ack => type_cast_1931_inst_req_0); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	228 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (5) 
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/word_access_start/$exit
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/word_access_start/word_0/$exit
      -- CP-element group 240: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Sample/word_access_start/word_0/ra
      -- 
    ra_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1911_load_0_ack_0, ack => zeropad3D_CP_2152_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	228 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	250 
    -- CP-element group 241:  members (9) 
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/word_access_complete/$exit
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/word_access_complete/word_0/$exit
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/word_access_complete/word_0/ca
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/ptr_deref_1911_Merge/$entry
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/ptr_deref_1911_Merge/$exit
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/ptr_deref_1911_Merge/merge_req
      -- CP-element group 241: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1911_Update/ptr_deref_1911_Merge/merge_ack
      -- 
    ca_5177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1911_load_0_ack_1, ack => zeropad3D_CP_2152_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	228 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (5) 
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/word_access_start/$exit
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/word_access_start/word_0/$exit
      -- CP-element group 242: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Sample/word_access_start/word_0/ra
      -- 
    ra_5216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1923_load_0_ack_0, ack => zeropad3D_CP_2152_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	228 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	250 
    -- CP-element group 243:  members (9) 
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/word_access_complete/$exit
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/word_access_complete/word_0/$exit
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/word_access_complete/word_0/ca
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/ptr_deref_1923_Merge/$entry
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/ptr_deref_1923_Merge/$exit
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/ptr_deref_1923_Merge/merge_req
      -- CP-element group 243: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/ptr_deref_1923_Update/ptr_deref_1923_Merge/merge_ack
      -- 
    ca_5227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1923_load_0_ack_1, ack => zeropad3D_CP_2152_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	237 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Sample/ra
      -- 
    ra_5241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1927_inst_ack_0, ack => zeropad3D_CP_2152_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	228 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	250 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1927_Update/ca
      -- 
    ca_5246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1927_inst_ack_1, ack => zeropad3D_CP_2152_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	239 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Sample/ra
      -- 
    ra_5255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1931_inst_ack_0, ack => zeropad3D_CP_2152_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	228 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	250 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1931_Update/ca
      -- 
    ca_5260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1931_inst_ack_1, ack => zeropad3D_CP_2152_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	235 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Sample/ra
      -- 
    ra_5269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1970_inst_ack_0, ack => zeropad3D_CP_2152_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	228 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/type_cast_1970_Update/ca
      -- 
    ca_5274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1970_inst_ack_1, ack => zeropad3D_CP_2152_elements(249)); -- 
    -- CP-element group 250:  join  fork  transition  place  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	233 
    -- CP-element group 250: 	241 
    -- CP-element group 250: 	243 
    -- CP-element group 250: 	245 
    -- CP-element group 250: 	247 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	920 
    -- CP-element group 250: 	921 
    -- CP-element group 250: 	922 
    -- CP-element group 250: 	923 
    -- CP-element group 250:  members (16) 
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460
      -- CP-element group 250: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012__exit__
      -- CP-element group 250: 	 branch_block_stmt_714/assign_stmt_1881_to_assign_stmt_2012/$exit
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2015/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2028/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Sample/rr
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Update/cr
      -- 
    rr_12320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(250), ack => type_cast_2025_inst_req_0); -- 
    cr_12325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(250), ack => type_cast_2025_inst_req_1); -- 
    zeropad3D_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(233) & zeropad3D_CP_2152_elements(241) & zeropad3D_CP_2152_elements(243) & zeropad3D_CP_2152_elements(245) & zeropad3D_CP_2152_elements(247) & zeropad3D_CP_2152_elements(249);
      gj_zeropad3D_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	930 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Sample/ra
      -- 
    ra_5286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2039_inst_ack_0, ack => zeropad3D_CP_2152_elements(251)); -- 
    -- CP-element group 252:  branch  transition  place  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	930 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (13) 
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048__entry__
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047__exit__
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/$exit
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Update/ca
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048_dead_link/$entry
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048_eval_test/$entry
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048_eval_test/$exit
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048_eval_test/branch_req
      -- CP-element group 252: 	 branch_block_stmt_714/R_cmp465_2049_place
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048_if_link/$entry
      -- CP-element group 252: 	 branch_block_stmt_714/if_stmt_2048_else_link/$entry
      -- 
    ca_5291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2039_inst_ack_1, ack => zeropad3D_CP_2152_elements(252)); -- 
    branch_req_5299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(252), ack => if_stmt_2048_branch_req_0); -- 
    -- CP-element group 253:  transition  place  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	931 
    -- CP-element group 253:  members (5) 
      -- CP-element group 253: 	 branch_block_stmt_714/if_stmt_2048_if_link/$exit
      -- CP-element group 253: 	 branch_block_stmt_714/if_stmt_2048_if_link/if_choice_transition
      -- CP-element group 253: 	 branch_block_stmt_714/whilex_xbody460_ifx_xthen496
      -- CP-element group 253: 	 branch_block_stmt_714/whilex_xbody460_ifx_xthen496_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_714/whilex_xbody460_ifx_xthen496_PhiReq/$exit
      -- 
    if_choice_transition_5304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2048_branch_ack_1, ack => zeropad3D_CP_2152_elements(253)); -- 
    -- CP-element group 254:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	258 
    -- CP-element group 254:  members (27) 
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079__entry__
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2054__exit__
      -- CP-element group 254: 	 branch_block_stmt_714/if_stmt_2048_else_link/$exit
      -- CP-element group 254: 	 branch_block_stmt_714/if_stmt_2048_else_link/else_choice_transition
      -- CP-element group 254: 	 branch_block_stmt_714/whilex_xbody460_lorx_xlhsx_xfalse467
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_update_start_
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_word_address_calculated
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_root_address_calculated
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/word_access_start/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/word_access_start/word_0/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/word_access_start/word_0/rr
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/word_access_complete/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/word_access_complete/word_0/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/word_access_complete/word_0/cr
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_update_start_
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Update/cr
      -- CP-element group 254: 	 branch_block_stmt_714/whilex_xbody460_lorx_xlhsx_xfalse467_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/whilex_xbody460_lorx_xlhsx_xfalse467_PhiReq/$exit
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2054_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2054_PhiAck/$entry
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2054_PhiAck/$exit
      -- CP-element group 254: 	 branch_block_stmt_714/merge_stmt_2054_PhiAck/dummy
      -- 
    else_choice_transition_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2048_branch_ack_0, ack => zeropad3D_CP_2152_elements(254)); -- 
    rr_5329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(254), ack => LOAD_row_high_2056_load_0_req_0); -- 
    cr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(254), ack => LOAD_row_high_2056_load_0_req_1); -- 
    cr_5359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(254), ack => type_cast_2060_inst_req_1); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (5) 
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/word_access_start/$exit
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/word_access_start/word_0/$exit
      -- CP-element group 255: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Sample/word_access_start/word_0/ra
      -- 
    ra_5330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2056_load_0_ack_0, ack => zeropad3D_CP_2152_elements(255)); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (12) 
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/word_access_complete/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/word_access_complete/word_0/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/word_access_complete/word_0/ca
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/LOAD_row_high_2056_Merge/$entry
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/LOAD_row_high_2056_Merge/$exit
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/LOAD_row_high_2056_Merge/merge_req
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/LOAD_row_high_2056_Update/LOAD_row_high_2056_Merge/merge_ack
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Sample/rr
      -- 
    ca_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2056_load_0_ack_1, ack => zeropad3D_CP_2152_elements(256)); -- 
    rr_5354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(256), ack => type_cast_2060_inst_req_0); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Sample/ra
      -- 
    ra_5355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2060_inst_ack_0, ack => zeropad3D_CP_2152_elements(257)); -- 
    -- CP-element group 258:  branch  transition  place  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	254 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (13) 
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080__entry__
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079__exit__
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/$exit
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_714/assign_stmt_2057_to_assign_stmt_2079/type_cast_2060_Update/ca
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080_dead_link/$entry
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080_eval_test/$entry
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080_eval_test/$exit
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080_eval_test/branch_req
      -- CP-element group 258: 	 branch_block_stmt_714/R_cmp476_2081_place
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080_if_link/$entry
      -- CP-element group 258: 	 branch_block_stmt_714/if_stmt_2080_else_link/$entry
      -- 
    ca_5360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2060_inst_ack_1, ack => zeropad3D_CP_2152_elements(258)); -- 
    branch_req_5368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(258), ack => if_stmt_2080_branch_req_0); -- 
    -- CP-element group 259:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	261 
    -- CP-element group 259: 	262 
    -- CP-element group 259:  members (18) 
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2086__exit__
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098__entry__
      -- CP-element group 259: 	 branch_block_stmt_714/if_stmt_2080_if_link/$exit
      -- CP-element group 259: 	 branch_block_stmt_714/if_stmt_2080_if_link/if_choice_transition
      -- CP-element group 259: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_lorx_xlhsx_xfalse478
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_update_start_
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_lorx_xlhsx_xfalse478_PhiReq/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_lorx_xlhsx_xfalse478_PhiReq/$exit
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2086_PhiReqMerge
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2086_PhiAck/$entry
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2086_PhiAck/$exit
      -- CP-element group 259: 	 branch_block_stmt_714/merge_stmt_2086_PhiAck/dummy
      -- 
    if_choice_transition_5373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2080_branch_ack_1, ack => zeropad3D_CP_2152_elements(259)); -- 
    rr_5390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => type_cast_2090_inst_req_0); -- 
    cr_5395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(259), ack => type_cast_2090_inst_req_1); -- 
    -- CP-element group 260:  transition  place  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	931 
    -- CP-element group 260:  members (5) 
      -- CP-element group 260: 	 branch_block_stmt_714/if_stmt_2080_else_link/$exit
      -- CP-element group 260: 	 branch_block_stmt_714/if_stmt_2080_else_link/else_choice_transition
      -- CP-element group 260: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_ifx_xthen496
      -- CP-element group 260: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_ifx_xthen496_PhiReq/$entry
      -- CP-element group 260: 	 branch_block_stmt_714/lorx_xlhsx_xfalse467_ifx_xthen496_PhiReq/$exit
      -- 
    else_choice_transition_5377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2080_branch_ack_0, ack => zeropad3D_CP_2152_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Sample/ra
      -- 
    ra_5391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2090_inst_ack_0, ack => zeropad3D_CP_2152_elements(261)); -- 
    -- CP-element group 262:  branch  transition  place  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	259 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (13) 
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098__exit__
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099__entry__
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/$exit
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_714/assign_stmt_2091_to_assign_stmt_2098/type_cast_2090_Update/ca
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099_dead_link/$entry
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099_eval_test/$entry
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099_eval_test/$exit
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099_eval_test/branch_req
      -- CP-element group 262: 	 branch_block_stmt_714/R_cmp483_2100_place
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099_if_link/$entry
      -- CP-element group 262: 	 branch_block_stmt_714/if_stmt_2099_else_link/$entry
      -- 
    ca_5396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2090_inst_ack_1, ack => zeropad3D_CP_2152_elements(262)); -- 
    branch_req_5404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(262), ack => if_stmt_2099_branch_req_0); -- 
    -- CP-element group 263:  transition  place  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	931 
    -- CP-element group 263:  members (5) 
      -- CP-element group 263: 	 branch_block_stmt_714/if_stmt_2099_if_link/$exit
      -- CP-element group 263: 	 branch_block_stmt_714/if_stmt_2099_if_link/if_choice_transition
      -- CP-element group 263: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_ifx_xthen496
      -- CP-element group 263: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_ifx_xthen496_PhiReq/$entry
      -- CP-element group 263: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_ifx_xthen496_PhiReq/$exit
      -- 
    if_choice_transition_5409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2099_branch_ack_1, ack => zeropad3D_CP_2152_elements(263)); -- 
    -- CP-element group 264:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264: 	266 
    -- CP-element group 264: 	268 
    -- CP-element group 264:  members (27) 
      -- CP-element group 264: 	 branch_block_stmt_714/merge_stmt_2105__exit__
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130__entry__
      -- CP-element group 264: 	 branch_block_stmt_714/if_stmt_2099_else_link/$exit
      -- CP-element group 264: 	 branch_block_stmt_714/if_stmt_2099_else_link/else_choice_transition
      -- CP-element group 264: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_lorx_xlhsx_xfalse485
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_update_start_
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_word_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_root_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/word_access_start/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/word_access_start/word_0/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/word_access_start/word_0/rr
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/word_access_complete/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/word_access_complete/word_0/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/word_access_complete/word_0/cr
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_update_start_
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Update/cr
      -- CP-element group 264: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_lorx_xlhsx_xfalse485_PhiReq/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/lorx_xlhsx_xfalse478_lorx_xlhsx_xfalse485_PhiReq/$exit
      -- CP-element group 264: 	 branch_block_stmt_714/merge_stmt_2105_PhiReqMerge
      -- CP-element group 264: 	 branch_block_stmt_714/merge_stmt_2105_PhiAck/$entry
      -- CP-element group 264: 	 branch_block_stmt_714/merge_stmt_2105_PhiAck/$exit
      -- CP-element group 264: 	 branch_block_stmt_714/merge_stmt_2105_PhiAck/dummy
      -- 
    else_choice_transition_5413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2099_branch_ack_0, ack => zeropad3D_CP_2152_elements(264)); -- 
    rr_5434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(264), ack => LOAD_col_high_2107_load_0_req_0); -- 
    cr_5445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(264), ack => LOAD_col_high_2107_load_0_req_1); -- 
    cr_5464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(264), ack => type_cast_2111_inst_req_1); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/word_access_start/$exit
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/word_access_start/word_0/$exit
      -- CP-element group 265: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Sample/word_access_start/word_0/ra
      -- 
    ra_5435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2107_load_0_ack_0, ack => zeropad3D_CP_2152_elements(265)); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (12) 
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/word_access_complete/$exit
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/word_access_complete/word_0/$exit
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/word_access_complete/word_0/ca
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/LOAD_col_high_2107_Merge/$entry
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/LOAD_col_high_2107_Merge/$exit
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/LOAD_col_high_2107_Merge/merge_req
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/LOAD_col_high_2107_Update/LOAD_col_high_2107_Merge/merge_ack
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Sample/rr
      -- 
    ca_5446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2107_load_0_ack_1, ack => zeropad3D_CP_2152_elements(266)); -- 
    rr_5459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(266), ack => type_cast_2111_inst_req_0); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Sample/ra
      -- 
    ra_5460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2111_inst_ack_0, ack => zeropad3D_CP_2152_elements(267)); -- 
    -- CP-element group 268:  branch  transition  place  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	264 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (13) 
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131__entry__
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130__exit__
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131_else_link/$entry
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/$exit
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_714/assign_stmt_2108_to_assign_stmt_2130/type_cast_2111_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131_dead_link/$entry
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131_eval_test/$entry
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131_eval_test/$exit
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131_eval_test/branch_req
      -- CP-element group 268: 	 branch_block_stmt_714/R_cmp494_2132_place
      -- CP-element group 268: 	 branch_block_stmt_714/if_stmt_2131_if_link/$entry
      -- 
    ca_5465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2111_inst_ack_1, ack => zeropad3D_CP_2152_elements(268)); -- 
    branch_req_5473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(268), ack => if_stmt_2131_branch_req_0); -- 
    -- CP-element group 269:  fork  transition  place  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	285 
    -- CP-element group 269: 	286 
    -- CP-element group 269: 	288 
    -- CP-element group 269: 	290 
    -- CP-element group 269: 	292 
    -- CP-element group 269: 	294 
    -- CP-element group 269: 	296 
    -- CP-element group 269: 	298 
    -- CP-element group 269: 	300 
    -- CP-element group 269: 	303 
    -- CP-element group 269:  members (46) 
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300__entry__
      -- CP-element group 269: 	 branch_block_stmt_714/merge_stmt_2195__exit__
      -- CP-element group 269: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xelse517
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Update/req
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Update/cr
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_update_start
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_complete/req
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Sample/rr
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Update/cr
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_update_start
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_complete/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/word_access_complete/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Update/req
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/word_access_complete/word_0/cr
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_complete/req
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_complete/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Update/cr
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/word_access_complete/word_0/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_update_start_
      -- CP-element group 269: 	 branch_block_stmt_714/if_stmt_2131_if_link/$exit
      -- CP-element group 269: 	 branch_block_stmt_714/if_stmt_2131_if_link/if_choice_transition
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/word_access_complete/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/word_access_complete/word_0/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/word_access_complete/word_0/cr
      -- CP-element group 269: 	 branch_block_stmt_714/merge_stmt_2195_PhiReqMerge
      -- CP-element group 269: 	 branch_block_stmt_714/merge_stmt_2195_PhiAck/dummy
      -- CP-element group 269: 	 branch_block_stmt_714/merge_stmt_2195_PhiAck/$exit
      -- CP-element group 269: 	 branch_block_stmt_714/merge_stmt_2195_PhiAck/$entry
      -- CP-element group 269: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xelse517_PhiReq/$exit
      -- CP-element group 269: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xelse517_PhiReq/$entry
      -- 
    if_choice_transition_5478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2131_branch_ack_1, ack => zeropad3D_CP_2152_elements(269)); -- 
    req_5686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => array_obj_ref_2269_index_offset_req_1); -- 
    cr_5641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => type_cast_2199_inst_req_1); -- 
    req_5811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => addr_of_2295_final_reg_req_1); -- 
    rr_5636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => type_cast_2199_inst_req_0); -- 
    cr_5765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => type_cast_2288_inst_req_1); -- 
    req_5796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => array_obj_ref_2294_index_offset_req_1); -- 
    cr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => ptr_deref_2274_load_0_req_1); -- 
    req_5701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => addr_of_2270_final_reg_req_1); -- 
    cr_5655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => type_cast_2263_inst_req_1); -- 
    cr_5861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(269), ack => ptr_deref_2298_store_0_req_1); -- 
    -- CP-element group 270:  transition  place  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	931 
    -- CP-element group 270:  members (5) 
      -- CP-element group 270: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xthen496
      -- CP-element group 270: 	 branch_block_stmt_714/if_stmt_2131_else_link/else_choice_transition
      -- CP-element group 270: 	 branch_block_stmt_714/if_stmt_2131_else_link/$exit
      -- CP-element group 270: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xthen496_PhiReq/$entry
      -- CP-element group 270: 	 branch_block_stmt_714/lorx_xlhsx_xfalse485_ifx_xthen496_PhiReq/$exit
      -- 
    else_choice_transition_5482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2131_branch_ack_0, ack => zeropad3D_CP_2152_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	931 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Sample/ra
      -- CP-element group 271: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_sample_completed_
      -- 
    ra_5496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_0, ack => zeropad3D_CP_2152_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	931 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	275 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Update/ca
      -- CP-element group 272: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Update/$exit
      -- 
    ca_5501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_1, ack => zeropad3D_CP_2152_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	931 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Sample/ra
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_sample_completed_
      -- 
    ra_5510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_0, ack => zeropad3D_CP_2152_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	931 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Update/ca
      -- CP-element group 274: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_update_completed_
      -- 
    ca_5515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_1, ack => zeropad3D_CP_2152_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	272 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Sample/rr
      -- CP-element group 275: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Sample/$entry
      -- 
    rr_5523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(275), ack => type_cast_2180_inst_req_0); -- 
    zeropad3D_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(272) & zeropad3D_CP_2152_elements(274);
      gj_zeropad3D_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Sample/ra
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_sample_completed_
      -- 
    ra_5524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_0, ack => zeropad3D_CP_2152_elements(276)); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	931 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (16) 
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_scale_1/$entry
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_resize_1/index_resize_ack
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_resize_1/index_resize_req
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_resize_1/$exit
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_resize_1/$entry
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_computed_1
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_scaled_1
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_resized_1
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Sample/req
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Update/ca
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_scale_1/scale_rename_ack
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_scale_1/scale_rename_req
      -- CP-element group 277: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_index_scale_1/$exit
      -- 
    ca_5529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_1, ack => zeropad3D_CP_2152_elements(277)); -- 
    req_5554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(277), ack => array_obj_ref_2186_index_offset_req_0); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	284 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Sample/ack
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_sample_complete
      -- 
    ack_5555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2186_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(278)); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	931 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (11) 
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_offset_calculated
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_root_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_request/req
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_request/$entry
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_base_plus_offset/sum_rename_ack
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_base_plus_offset/sum_rename_req
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_base_plus_offset/$exit
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_base_plus_offset/$entry
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Update/ack
      -- CP-element group 279: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Update/$exit
      -- 
    ack_5560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2186_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(279)); -- 
    req_5569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(279), ack => addr_of_2187_final_reg_req_0); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_request/ack
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_request/$exit
      -- 
    ack_5570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2187_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(280)); -- 
    -- CP-element group 281:  join  fork  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	931 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (28) 
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/word_access_start/word_0/rr
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/word_access_start/word_0/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/word_access_start/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/ptr_deref_2190_Split/split_ack
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/ptr_deref_2190_Split/split_req
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/ptr_deref_2190_Split/$exit
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/ptr_deref_2190_Split/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_word_addrgen/root_register_ack
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_word_addrgen/root_register_req
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_word_addrgen/$exit
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_word_addrgen/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_plus_offset/sum_rename_ack
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_plus_offset/sum_rename_req
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_plus_offset/$exit
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_plus_offset/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_addr_resize/base_resize_ack
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_addr_resize/base_resize_req
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_addr_resize/$exit
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_addr_resize/$entry
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_address_resized
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_root_address_calculated
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_word_address_calculated
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_base_address_calculated
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_update_completed_
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_complete/ack
      -- CP-element group 281: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_complete/$exit
      -- 
    ack_5575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2187_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(281)); -- 
    rr_5613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(281), ack => ptr_deref_2190_store_0_req_0); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (5) 
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/word_access_start/word_0/ra
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/word_access_start/word_0/$exit
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/word_access_start/$exit
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_sample_completed_
      -- 
    ra_5614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2190_store_0_ack_0, ack => zeropad3D_CP_2152_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	931 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (5) 
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/word_access_complete/$exit
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/word_access_complete/word_0/ca
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/word_access_complete/word_0/$exit
      -- 
    ca_5625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2190_store_0_ack_1, ack => zeropad3D_CP_2152_elements(283)); -- 
    -- CP-element group 284:  join  transition  place  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: 	278 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	932 
    -- CP-element group 284:  members (5) 
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193__exit__
      -- CP-element group 284: 	 branch_block_stmt_714/ifx_xthen496_ifx_xend565
      -- CP-element group 284: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/$exit
      -- CP-element group 284: 	 branch_block_stmt_714/ifx_xthen496_ifx_xend565_PhiReq/$exit
      -- CP-element group 284: 	 branch_block_stmt_714/ifx_xthen496_ifx_xend565_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(283) & zeropad3D_CP_2152_elements(278);
      gj_zeropad3D_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	269 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Sample/ra
      -- CP-element group 285: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_sample_completed_
      -- 
    ra_5637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => zeropad3D_CP_2152_elements(285)); -- 
    -- CP-element group 286:  fork  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	269 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286: 	295 
    -- CP-element group 286:  members (9) 
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_Update/ca
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Sample/rr
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2199_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Sample/rr
      -- CP-element group 286: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Sample/$entry
      -- 
    ca_5642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => zeropad3D_CP_2152_elements(286)); -- 
    rr_5650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(286), ack => type_cast_2263_inst_req_0); -- 
    rr_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(286), ack => type_cast_2288_inst_req_0); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Sample/ra
      -- CP-element group 287: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Sample/$exit
      -- 
    ra_5651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2263_inst_ack_0, ack => zeropad3D_CP_2152_elements(287)); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	269 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (16) 
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_scale_1/scale_rename_ack
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_scale_1/scale_rename_req
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_scale_1/$exit
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_scale_1/$entry
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_resize_1/index_resize_ack
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_resize_1/index_resize_req
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_resize_1/$exit
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_resize_1/$entry
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_computed_1
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_scaled_1
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_index_resized_1
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Update/ca
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2263_update_completed_
      -- 
    ca_5656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2263_inst_ack_1, ack => zeropad3D_CP_2152_elements(288)); -- 
    req_5681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(288), ack => array_obj_ref_2269_index_offset_req_0); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	304 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_sample_complete
      -- 
    ack_5682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2269_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(289)); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	269 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (11) 
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_base_plus_offset/$entry
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_base_plus_offset/$exit
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_base_plus_offset/sum_rename_req
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_base_plus_offset/sum_rename_ack
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_request/$entry
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_final_index_sum_regn_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_offset_calculated
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2269_root_address_calculated
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_request/req
      -- 
    ack_5687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2269_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(290)); -- 
    req_5696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(290), ack => addr_of_2270_final_reg_req_0); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_request/ack
      -- CP-element group 291: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_request/$exit
      -- 
    ack_5697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2270_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(291)); -- 
    -- CP-element group 292:  join  fork  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	269 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (24) 
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/word_access_start/$entry
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/word_access_start/word_0/$entry
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_word_addrgen/root_register_ack
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_word_addrgen/root_register_req
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_word_addrgen/$exit
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_word_addrgen/$entry
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_plus_offset/sum_rename_ack
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_plus_offset/sum_rename_req
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_plus_offset/$exit
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_plus_offset/$entry
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_addr_resize/base_resize_ack
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_addr_resize/base_resize_req
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_addr_resize/$exit
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/word_access_start/word_0/rr
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_addr_resize/$entry
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_address_resized
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_root_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_word_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_base_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_complete/ack
      -- CP-element group 292: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2270_complete/$exit
      -- 
    ack_5702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2270_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(292)); -- 
    rr_5735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(292), ack => ptr_deref_2274_load_0_req_0); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293:  members (5) 
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/word_access_start/$exit
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/word_access_start/word_0/ra
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Sample/word_access_start/word_0/$exit
      -- CP-element group 293: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_sample_completed_
      -- 
    ra_5736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2274_load_0_ack_0, ack => zeropad3D_CP_2152_elements(293)); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	269 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	301 
    -- CP-element group 294:  members (9) 
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/ptr_deref_2274_Merge/merge_ack
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/ptr_deref_2274_Merge/merge_req
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/ptr_deref_2274_Merge/$exit
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/ptr_deref_2274_Merge/$entry
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/word_access_complete/word_0/ca
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/word_access_complete/word_0/$exit
      -- CP-element group 294: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2274_Update/word_access_complete/$exit
      -- 
    ca_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2274_load_0_ack_1, ack => zeropad3D_CP_2152_elements(294)); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	286 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Sample/ra
      -- CP-element group 295: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_sample_completed_
      -- 
    ra_5761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_0, ack => zeropad3D_CP_2152_elements(295)); -- 
    -- CP-element group 296:  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	269 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (16) 
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_resized_1
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_scaled_1
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Update/ca
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_scale_1/scale_rename_ack
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/type_cast_2288_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_scale_1/scale_rename_req
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_scale_1/$exit
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_scale_1/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_resize_1/index_resize_ack
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Sample/req
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_resize_1/index_resize_req
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_resize_1/$exit
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_resize_1/$entry
      -- CP-element group 296: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_index_computed_1
      -- 
    ca_5766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_1, ack => zeropad3D_CP_2152_elements(296)); -- 
    req_5791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(296), ack => array_obj_ref_2294_index_offset_req_0); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	304 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_sample_complete
      -- CP-element group 297: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Sample/ack
      -- 
    ack_5792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2294_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(297)); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	269 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (11) 
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_offset_calculated
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_root_address_calculated
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_request/req
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_base_plus_offset/sum_rename_ack
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_base_plus_offset/sum_rename_req
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_base_plus_offset/$exit
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_base_plus_offset/$entry
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/array_obj_ref_2294_final_index_sum_regn_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_request/$entry
      -- 
    ack_5797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2294_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(298)); -- 
    req_5806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(298), ack => addr_of_2295_final_reg_req_0); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_request/ack
      -- CP-element group 299: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_request/$exit
      -- 
    ack_5807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2295_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	269 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (19) 
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_complete/ack
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_addr_resize/base_resize_ack
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_address_resized
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_word_addrgen/$entry
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_addr_resize/base_resize_req
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/addr_of_2295_complete/$exit
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_addr_resize/$exit
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_root_address_calculated
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_plus_offset/sum_rename_ack
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_addr_resize/$entry
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_word_address_calculated
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_address_calculated
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_plus_offset/sum_rename_req
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_plus_offset/$entry
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_base_plus_offset/$exit
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_word_addrgen/$exit
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_word_addrgen/root_register_req
      -- CP-element group 300: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_word_addrgen/root_register_ack
      -- 
    ack_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2295_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	294 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (9) 
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/ptr_deref_2298_Split/$entry
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/ptr_deref_2298_Split/$exit
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/ptr_deref_2298_Split/split_req
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/ptr_deref_2298_Split/split_ack
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/word_access_start/$entry
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/word_access_start/word_0/$entry
      -- CP-element group 301: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/word_access_start/word_0/rr
      -- 
    rr_5850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(301), ack => ptr_deref_2298_store_0_req_0); -- 
    zeropad3D_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(294) & zeropad3D_CP_2152_elements(300);
      gj_zeropad3D_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (5) 
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_sample_completed_
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/word_access_start/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/word_access_start/word_0/$exit
      -- CP-element group 302: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Sample/word_access_start/word_0/ra
      -- 
    ra_5851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2298_store_0_ack_0, ack => zeropad3D_CP_2152_elements(302)); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	269 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (5) 
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_update_completed_
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/$exit
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/word_access_complete/$exit
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/word_access_complete/word_0/$exit
      -- CP-element group 303: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/ptr_deref_2298_Update/word_access_complete/word_0/ca
      -- 
    ca_5862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2298_store_0_ack_1, ack => zeropad3D_CP_2152_elements(303)); -- 
    -- CP-element group 304:  join  transition  place  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	289 
    -- CP-element group 304: 	297 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	932 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300__exit__
      -- CP-element group 304: 	 branch_block_stmt_714/ifx_xelse517_ifx_xend565
      -- CP-element group 304: 	 branch_block_stmt_714/assign_stmt_2200_to_assign_stmt_2300/$exit
      -- CP-element group 304: 	 branch_block_stmt_714/ifx_xelse517_ifx_xend565_PhiReq/$entry
      -- CP-element group 304: 	 branch_block_stmt_714/ifx_xelse517_ifx_xend565_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(289) & zeropad3D_CP_2152_elements(297) & zeropad3D_CP_2152_elements(303);
      gj_zeropad3D_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	932 
    -- CP-element group 305: successors 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Sample/ra
      -- 
    ra_5874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_0, ack => zeropad3D_CP_2152_elements(305)); -- 
    -- CP-element group 306:  branch  transition  place  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	932 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (13) 
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321__entry__
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320__exit__
      -- CP-element group 306: 	 branch_block_stmt_714/R_cmp573_2322_place
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/$exit
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Update/ca
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321_dead_link/$entry
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321_eval_test/$entry
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321_eval_test/$exit
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321_eval_test/branch_req
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321_if_link/$entry
      -- CP-element group 306: 	 branch_block_stmt_714/if_stmt_2321_else_link/$entry
      -- 
    ca_5879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_1, ack => zeropad3D_CP_2152_elements(306)); -- 
    branch_req_5887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(306), ack => if_stmt_2321_branch_req_0); -- 
    -- CP-element group 307:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	941 
    -- CP-element group 307: 	942 
    -- CP-element group 307: 	944 
    -- CP-element group 307: 	945 
    -- CP-element group 307: 	947 
    -- CP-element group 307: 	948 
    -- CP-element group 307:  members (40) 
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2333__exit__
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2333__entry__
      -- CP-element group 307: 	 branch_block_stmt_714/merge_stmt_2327__exit__
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xend565_ifx_xthen575
      -- CP-element group 307: 	 branch_block_stmt_714/if_stmt_2321_if_link/$exit
      -- CP-element group 307: 	 branch_block_stmt_714/if_stmt_2321_if_link/if_choice_transition
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2333/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/assign_stmt_2333/$exit
      -- CP-element group 307: 	 branch_block_stmt_714/merge_stmt_2327_PhiReqMerge
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/cr
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/rr
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Update/cr
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/merge_stmt_2327_PhiAck/dummy
      -- CP-element group 307: 	 branch_block_stmt_714/merge_stmt_2327_PhiAck/$exit
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/merge_stmt_2327_PhiAck/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xend565_ifx_xthen575_PhiReq/$exit
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xend565_ifx_xthen575_PhiReq/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Update/cr
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Sample/rr
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Sample/rr
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Sample/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Sample/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/$entry
      -- CP-element group 307: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/$entry
      -- 
    if_choice_transition_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2321_branch_ack_1, ack => zeropad3D_CP_2152_elements(307)); -- 
    cr_12561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2437_inst_req_1); -- 
    rr_12556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2437_inst_req_0); -- 
    cr_12515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2424_inst_req_1); -- 
    cr_12538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2431_inst_req_1); -- 
    rr_12510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2424_inst_req_0); -- 
    rr_12533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(307), ack => type_cast_2431_inst_req_0); -- 
    -- CP-element group 308:  fork  transition  place  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308: 	310 
    -- CP-element group 308: 	311 
    -- CP-element group 308: 	312 
    -- CP-element group 308: 	314 
    -- CP-element group 308: 	317 
    -- CP-element group 308: 	319 
    -- CP-element group 308: 	320 
    -- CP-element group 308: 	321 
    -- CP-element group 308: 	323 
    -- CP-element group 308:  members (54) 
      -- CP-element group 308: 	 branch_block_stmt_714/merge_stmt_2335__exit__
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413__entry__
      -- CP-element group 308: 	 branch_block_stmt_714/ifx_xend565_ifx_xelse580
      -- CP-element group 308: 	 branch_block_stmt_714/if_stmt_2321_else_link/$exit
      -- CP-element group 308: 	 branch_block_stmt_714/if_stmt_2321_else_link/else_choice_transition
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Sample/rr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/word_access_start/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/word_access_start/word_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/word_access_start/word_0/rr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/word_access_complete/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/word_access_complete/word_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/word_access_complete/word_0/cr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_word_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_root_address_calculated
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/word_access_start/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/word_access_start/word_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/word_access_start/word_0/rr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/word_access_complete/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/word_access_complete/word_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/word_access_complete/word_0/cr
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_update_start_
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Update/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Update/cr
      -- CP-element group 308: 	 branch_block_stmt_714/merge_stmt_2335_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_714/merge_stmt_2335_PhiAck/dummy
      -- CP-element group 308: 	 branch_block_stmt_714/merge_stmt_2335_PhiAck/$exit
      -- CP-element group 308: 	 branch_block_stmt_714/merge_stmt_2335_PhiAck/$entry
      -- CP-element group 308: 	 branch_block_stmt_714/ifx_xend565_ifx_xelse580_PhiReq/$exit
      -- CP-element group 308: 	 branch_block_stmt_714/ifx_xend565_ifx_xelse580_PhiReq/$entry
      -- 
    else_choice_transition_5896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2321_branch_ack_0, ack => zeropad3D_CP_2152_elements(308)); -- 
    rr_5912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => type_cast_2345_inst_req_0); -- 
    cr_5917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => type_cast_2345_inst_req_1); -- 
    rr_5934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => LOAD_col_high_2348_load_0_req_0); -- 
    cr_5945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => LOAD_col_high_2348_load_0_req_1); -- 
    cr_5964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => type_cast_2352_inst_req_1); -- 
    cr_5978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => type_cast_2372_inst_req_1); -- 
    cr_5992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => type_cast_2389_inst_req_1); -- 
    rr_6009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => LOAD_row_high_2392_load_0_req_0); -- 
    cr_6020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => LOAD_row_high_2392_load_0_req_1); -- 
    cr_6039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(308), ack => type_cast_2396_inst_req_1); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Sample/ra
      -- 
    ra_5913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2345_inst_ack_0, ack => zeropad3D_CP_2152_elements(309)); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	315 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2345_Update/ca
      -- 
    ca_5918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2345_inst_ack_1, ack => zeropad3D_CP_2152_elements(310)); -- 
    -- CP-element group 311:  transition  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	308 
    -- CP-element group 311: successors 
    -- CP-element group 311:  members (5) 
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/word_access_start/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/word_access_start/word_0/$exit
      -- CP-element group 311: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Sample/word_access_start/word_0/ra
      -- 
    ra_5935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2348_load_0_ack_0, ack => zeropad3D_CP_2152_elements(311)); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	308 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (12) 
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/word_access_complete/$exit
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/word_access_complete/word_0/$exit
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/word_access_complete/word_0/ca
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/LOAD_col_high_2348_Merge/$entry
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/LOAD_col_high_2348_Merge/$exit
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/LOAD_col_high_2348_Merge/merge_req
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_col_high_2348_Update/LOAD_col_high_2348_Merge/merge_ack
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Sample/rr
      -- 
    ca_5946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2348_load_0_ack_1, ack => zeropad3D_CP_2152_elements(312)); -- 
    rr_5959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(312), ack => type_cast_2352_inst_req_0); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Sample/ra
      -- 
    ra_5960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_0, ack => zeropad3D_CP_2152_elements(313)); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	308 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2352_Update/ca
      -- 
    ca_5965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_1, ack => zeropad3D_CP_2152_elements(314)); -- 
    -- CP-element group 315:  join  transition  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	310 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_sample_start_
      -- CP-element group 315: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Sample/rr
      -- 
    rr_5973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(315), ack => type_cast_2372_inst_req_0); -- 
    zeropad3D_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(310) & zeropad3D_CP_2152_elements(314);
      gj_zeropad3D_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_sample_completed_
      -- CP-element group 316: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Sample/ra
      -- 
    ra_5974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2372_inst_ack_0, ack => zeropad3D_CP_2152_elements(316)); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	308 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2372_Update/ca
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Sample/rr
      -- 
    ca_5979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2372_inst_ack_1, ack => zeropad3D_CP_2152_elements(317)); -- 
    rr_5987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(317), ack => type_cast_2389_inst_req_0); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Sample/ra
      -- 
    ra_5988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_0, ack => zeropad3D_CP_2152_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	308 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	324 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2389_Update/ca
      -- 
    ca_5993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2389_inst_ack_1, ack => zeropad3D_CP_2152_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	308 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (5) 
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/word_access_start/$exit
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/word_access_start/word_0/$exit
      -- CP-element group 320: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Sample/word_access_start/word_0/ra
      -- 
    ra_6010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2392_load_0_ack_0, ack => zeropad3D_CP_2152_elements(320)); -- 
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	308 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (12) 
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/word_access_complete/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/word_access_complete/word_0/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/word_access_complete/word_0/ca
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/LOAD_row_high_2392_Merge/$entry
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/LOAD_row_high_2392_Merge/$exit
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/LOAD_row_high_2392_Merge/merge_req
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/LOAD_row_high_2392_Update/LOAD_row_high_2392_Merge/merge_ack
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_sample_start_
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Sample/rr
      -- 
    ca_6021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2392_load_0_ack_1, ack => zeropad3D_CP_2152_elements(321)); -- 
    rr_6034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(321), ack => type_cast_2396_inst_req_0); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_sample_completed_
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Sample/ra
      -- 
    ra_6035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2396_inst_ack_0, ack => zeropad3D_CP_2152_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	308 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_update_completed_
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Update/$exit
      -- CP-element group 323: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/type_cast_2396_Update/ca
      -- 
    ca_6040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2396_inst_ack_1, ack => zeropad3D_CP_2152_elements(323)); -- 
    -- CP-element group 324:  branch  join  transition  place  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	319 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (10) 
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413__exit__
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414__entry__
      -- CP-element group 324: 	 branch_block_stmt_714/assign_stmt_2341_to_assign_stmt_2413/$exit
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414_dead_link/$entry
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414_eval_test/$entry
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414_eval_test/$exit
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414_eval_test/branch_req
      -- CP-element group 324: 	 branch_block_stmt_714/R_cmp608_2415_place
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414_if_link/$entry
      -- CP-element group 324: 	 branch_block_stmt_714/if_stmt_2414_else_link/$entry
      -- 
    branch_req_6048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(324), ack => if_stmt_2414_branch_req_0); -- 
    zeropad3D_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(319) & zeropad3D_CP_2152_elements(323);
      gj_zeropad3D_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: 	328 
    -- CP-element group 325: 	330 
    -- CP-element group 325: 	331 
    -- CP-element group 325: 	332 
    -- CP-element group 325: 	334 
    -- CP-element group 325: 	335 
    -- CP-element group 325: 	336 
    -- CP-element group 325: 	337 
    -- CP-element group 325: 	338 
    -- CP-element group 325: 	339 
    -- CP-element group 325: 	340 
    -- CP-element group 325: 	341 
    -- CP-element group 325: 	342 
    -- CP-element group 325: 	344 
    -- CP-element group 325: 	346 
    -- CP-element group 325: 	348 
    -- CP-element group 325:  members (127) 
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587__entry__
      -- CP-element group 325: 	 branch_block_stmt_714/merge_stmt_2442__exit__
      -- CP-element group 325: 	 branch_block_stmt_714/if_stmt_2414_if_link/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/if_stmt_2414_if_link/if_choice_transition
      -- CP-element group 325: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_word_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_root_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/word_access_start/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/word_access_start/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/word_access_start/word_0/rr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/word_access_complete/word_0/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Update/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_word_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_root_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/word_access_start/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/word_access_start/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/word_access_start/word_0/rr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/word_access_complete/word_0/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Update/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_word_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_root_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/word_access_start/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/word_access_start/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/word_access_start/word_0/rr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/word_access_complete/word_0/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_word_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_root_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/word_access_start/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/word_access_start/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/word_access_start/word_0/rr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/word_access_complete/word_0/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_word_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_root_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_address_resized
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_addr_resize/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_addr_resize/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_addr_resize/base_resize_req
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_addr_resize/base_resize_ack
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_plus_offset/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_plus_offset/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_plus_offset/sum_rename_req
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_base_plus_offset/sum_rename_ack
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_word_addrgen/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_word_addrgen/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_word_addrgen/root_register_req
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_word_addrgen/root_register_ack
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/word_access_start/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/word_access_start/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/word_access_start/word_0/rr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/word_access_complete/word_0/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_word_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_root_address_calculated
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_address_resized
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_addr_resize/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_addr_resize/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_addr_resize/base_resize_req
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_addr_resize/base_resize_ack
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_plus_offset/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_plus_offset/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_plus_offset/sum_rename_req
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_base_plus_offset/sum_rename_ack
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_word_addrgen/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_word_addrgen/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_word_addrgen/root_register_req
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_word_addrgen/root_register_ack
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/word_access_start/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/word_access_start/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/word_access_start/word_0/rr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/word_access_complete/word_0/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Update/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Update/cr
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_update_start_
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Update/cr
      -- CP-element group 325: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/ifx_xelse580_whilex_xend618_PhiReq/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/merge_stmt_2442_PhiAck/dummy
      -- CP-element group 325: 	 branch_block_stmt_714/merge_stmt_2442_PhiAck/$exit
      -- CP-element group 325: 	 branch_block_stmt_714/merge_stmt_2442_PhiAck/$entry
      -- CP-element group 325: 	 branch_block_stmt_714/merge_stmt_2442_PhiReqMerge
      -- 
    if_choice_transition_6053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2414_branch_ack_1, ack => zeropad3D_CP_2152_elements(325)); -- 
    rr_6078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_col_high_2445_load_0_req_0); -- 
    cr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_col_high_2445_load_0_req_1); -- 
    cr_6108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => type_cast_2449_inst_req_1); -- 
    rr_6125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_row_high_2458_load_0_req_0); -- 
    cr_6136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_row_high_2458_load_0_req_1); -- 
    cr_6155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => type_cast_2462_inst_req_1); -- 
    rr_6172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_pad_2471_load_0_req_0); -- 
    cr_6183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_pad_2471_load_0_req_1); -- 
    rr_6205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_depth_high_2474_load_0_req_0); -- 
    cr_6216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => LOAD_depth_high_2474_load_0_req_1); -- 
    rr_6255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => ptr_deref_2486_load_0_req_0); -- 
    cr_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => ptr_deref_2486_load_0_req_1); -- 
    rr_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => ptr_deref_2498_load_0_req_0); -- 
    cr_6316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => ptr_deref_2498_load_0_req_1); -- 
    cr_6335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => type_cast_2502_inst_req_1); -- 
    cr_6349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => type_cast_2506_inst_req_1); -- 
    cr_6363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(325), ack => type_cast_2545_inst_req_1); -- 
    -- CP-element group 326:  fork  transition  place  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	933 
    -- CP-element group 326: 	934 
    -- CP-element group 326: 	935 
    -- CP-element group 326: 	937 
    -- CP-element group 326: 	938 
    -- CP-element group 326:  members (22) 
      -- CP-element group 326: 	 branch_block_stmt_714/if_stmt_2414_else_link/$exit
      -- CP-element group 326: 	 branch_block_stmt_714/if_stmt_2414_else_link/else_choice_transition
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Update/cr
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2421/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/$entry
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Update/cr
      -- CP-element group 326: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/$entry
      -- 
    else_choice_transition_6057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2414_branch_ack_0, ack => zeropad3D_CP_2152_elements(326)); -- 
    rr_12461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(326), ack => type_cast_2433_inst_req_0); -- 
    cr_12489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(326), ack => type_cast_2439_inst_req_1); -- 
    rr_12484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(326), ack => type_cast_2439_inst_req_0); -- 
    cr_12466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(326), ack => type_cast_2433_inst_req_1); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/word_access_start/$exit
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/word_access_start/word_0/$exit
      -- CP-element group 327: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Sample/word_access_start/word_0/ra
      -- 
    ra_6079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2445_load_0_ack_0, ack => zeropad3D_CP_2152_elements(327)); -- 
    -- CP-element group 328:  fork  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	325 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328: 	345 
    -- CP-element group 328:  members (15) 
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/word_access_complete/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/word_access_complete/word_0/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/word_access_complete/word_0/ca
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/LOAD_col_high_2445_Merge/$entry
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/LOAD_col_high_2445_Merge/$exit
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/LOAD_col_high_2445_Merge/merge_req
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_col_high_2445_Update/LOAD_col_high_2445_Merge/merge_ack
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Sample/rr
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Sample/rr
      -- 
    ca_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2445_load_0_ack_1, ack => zeropad3D_CP_2152_elements(328)); -- 
    rr_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(328), ack => type_cast_2449_inst_req_0); -- 
    rr_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(328), ack => type_cast_2506_inst_req_0); -- 
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Sample/ra
      -- 
    ra_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2449_inst_ack_0, ack => zeropad3D_CP_2152_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	325 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	349 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2449_Update/ca
      -- 
    ca_6109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2449_inst_ack_1, ack => zeropad3D_CP_2152_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	325 
    -- CP-element group 331: successors 
    -- CP-element group 331:  members (5) 
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/word_access_start/$exit
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/word_access_start/word_0/$exit
      -- CP-element group 331: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Sample/word_access_start/word_0/ra
      -- 
    ra_6126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2458_load_0_ack_0, ack => zeropad3D_CP_2152_elements(331)); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	325 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (12) 
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/word_access_complete/$exit
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/word_access_complete/word_0/$exit
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/word_access_complete/word_0/ca
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/LOAD_row_high_2458_Merge/$entry
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/LOAD_row_high_2458_Merge/$exit
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/LOAD_row_high_2458_Merge/merge_req
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_row_high_2458_Update/LOAD_row_high_2458_Merge/merge_ack
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Sample/rr
      -- 
    ca_6137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2458_load_0_ack_1, ack => zeropad3D_CP_2152_elements(332)); -- 
    rr_6150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(332), ack => type_cast_2462_inst_req_0); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Sample/ra
      -- 
    ra_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2462_inst_ack_0, ack => zeropad3D_CP_2152_elements(333)); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	325 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	349 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2462_Update/ca
      -- 
    ca_6156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2462_inst_ack_1, ack => zeropad3D_CP_2152_elements(334)); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	325 
    -- CP-element group 335: successors 
    -- CP-element group 335:  members (5) 
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/word_access_start/$exit
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/word_access_start/word_0/$exit
      -- CP-element group 335: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Sample/word_access_start/word_0/ra
      -- 
    ra_6173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2471_load_0_ack_0, ack => zeropad3D_CP_2152_elements(335)); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	325 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	347 
    -- CP-element group 336:  members (12) 
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/word_access_complete/$exit
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/word_access_complete/word_0/$exit
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/word_access_complete/word_0/ca
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/LOAD_pad_2471_Merge/$entry
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/LOAD_pad_2471_Merge/$exit
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/LOAD_pad_2471_Merge/merge_req
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_pad_2471_Update/LOAD_pad_2471_Merge/merge_ack
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Sample/rr
      -- 
    ca_6184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2471_load_0_ack_1, ack => zeropad3D_CP_2152_elements(336)); -- 
    rr_6358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(336), ack => type_cast_2545_inst_req_0); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	325 
    -- CP-element group 337: successors 
    -- CP-element group 337:  members (5) 
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/word_access_start/$exit
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/word_access_start/word_0/$exit
      -- CP-element group 337: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Sample/word_access_start/word_0/ra
      -- 
    ra_6206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2474_load_0_ack_0, ack => zeropad3D_CP_2152_elements(337)); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	325 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	343 
    -- CP-element group 338:  members (12) 
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/word_access_complete/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/word_access_complete/word_0/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/word_access_complete/word_0/ca
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/LOAD_depth_high_2474_Merge/$entry
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/LOAD_depth_high_2474_Merge/$exit
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/LOAD_depth_high_2474_Merge/merge_req
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/LOAD_depth_high_2474_Update/LOAD_depth_high_2474_Merge/merge_ack
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Sample/rr
      -- 
    ca_6217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_2474_load_0_ack_1, ack => zeropad3D_CP_2152_elements(338)); -- 
    rr_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(338), ack => type_cast_2502_inst_req_0); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	325 
    -- CP-element group 339: successors 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/word_access_start/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/word_access_start/word_0/$exit
      -- CP-element group 339: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Sample/word_access_start/word_0/ra
      -- 
    ra_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2486_load_0_ack_0, ack => zeropad3D_CP_2152_elements(339)); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	325 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	349 
    -- CP-element group 340:  members (9) 
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/word_access_complete/$exit
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/word_access_complete/word_0/$exit
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/word_access_complete/word_0/ca
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/ptr_deref_2486_Merge/$entry
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/ptr_deref_2486_Merge/$exit
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/ptr_deref_2486_Merge/merge_req
      -- CP-element group 340: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2486_Update/ptr_deref_2486_Merge/merge_ack
      -- 
    ca_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2486_load_0_ack_1, ack => zeropad3D_CP_2152_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	325 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (5) 
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/word_access_start/$exit
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/word_access_start/word_0/$exit
      -- CP-element group 341: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Sample/word_access_start/word_0/ra
      -- 
    ra_6306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2498_load_0_ack_0, ack => zeropad3D_CP_2152_elements(341)); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	325 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	349 
    -- CP-element group 342:  members (9) 
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/word_access_complete/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/word_access_complete/word_0/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/word_access_complete/word_0/ca
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/ptr_deref_2498_Merge/$entry
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/ptr_deref_2498_Merge/$exit
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/ptr_deref_2498_Merge/merge_req
      -- CP-element group 342: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/ptr_deref_2498_Update/ptr_deref_2498_Merge/merge_ack
      -- 
    ca_6317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2498_load_0_ack_1, ack => zeropad3D_CP_2152_elements(342)); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	338 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Sample/ra
      -- 
    ra_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2502_inst_ack_0, ack => zeropad3D_CP_2152_elements(343)); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	325 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	349 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2502_Update/ca
      -- 
    ca_6336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2502_inst_ack_1, ack => zeropad3D_CP_2152_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	328 
    -- CP-element group 345: successors 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Sample/ra
      -- 
    ra_6345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_0, ack => zeropad3D_CP_2152_elements(345)); -- 
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	325 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	349 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2506_Update/ca
      -- 
    ca_6350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_1, ack => zeropad3D_CP_2152_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	336 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Sample/ra
      -- 
    ra_6359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2545_inst_ack_0, ack => zeropad3D_CP_2152_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	325 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/type_cast_2545_Update/ca
      -- 
    ca_6364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2545_inst_ack_1, ack => zeropad3D_CP_2152_elements(348)); -- 
    -- CP-element group 349:  join  fork  transition  place  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	330 
    -- CP-element group 349: 	334 
    -- CP-element group 349: 	340 
    -- CP-element group 349: 	342 
    -- CP-element group 349: 	344 
    -- CP-element group 349: 	346 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	966 
    -- CP-element group 349: 	967 
    -- CP-element group 349: 	968 
    -- CP-element group 349: 	970 
    -- CP-element group 349: 	971 
    -- CP-element group 349:  members (22) 
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587__exit__
      -- CP-element group 349: 	 branch_block_stmt_714/assign_stmt_2446_to_assign_stmt_2587/$exit
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2590/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Sample/rr
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Update/cr
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Sample/rr
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Update/cr
      -- 
    rr_12677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(349), ack => type_cast_2600_inst_req_0); -- 
    cr_12682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(349), ack => type_cast_2600_inst_req_1); -- 
    rr_12700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(349), ack => type_cast_2606_inst_req_0); -- 
    cr_12705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(349), ack => type_cast_2606_inst_req_1); -- 
    zeropad3D_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(330) & zeropad3D_CP_2152_elements(334) & zeropad3D_CP_2152_elements(340) & zeropad3D_CP_2152_elements(342) & zeropad3D_CP_2152_elements(344) & zeropad3D_CP_2152_elements(346) & zeropad3D_CP_2152_elements(348);
      gj_zeropad3D_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	978 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Sample/ra
      -- 
    ra_6376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2613_inst_ack_0, ack => zeropad3D_CP_2152_elements(350)); -- 
    -- CP-element group 351:  branch  transition  place  input  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	978 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (13) 
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622__entry__
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621__exit__
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/$exit
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Update/ca
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622_dead_link/$entry
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622_eval_test/$entry
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622_eval_test/$exit
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622_eval_test/branch_req
      -- CP-element group 351: 	 branch_block_stmt_714/R_cmp687_2623_place
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622_if_link/$entry
      -- CP-element group 351: 	 branch_block_stmt_714/if_stmt_2622_else_link/$entry
      -- 
    ca_6381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2613_inst_ack_1, ack => zeropad3D_CP_2152_elements(351)); -- 
    branch_req_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(351), ack => if_stmt_2622_branch_req_0); -- 
    -- CP-element group 352:  transition  place  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	979 
    -- CP-element group 352:  members (5) 
      -- CP-element group 352: 	 branch_block_stmt_714/if_stmt_2622_if_link/$exit
      -- CP-element group 352: 	 branch_block_stmt_714/if_stmt_2622_if_link/if_choice_transition
      -- CP-element group 352: 	 branch_block_stmt_714/whilex_xbody682_ifx_xthen717
      -- CP-element group 352: 	 branch_block_stmt_714/whilex_xbody682_ifx_xthen717_PhiReq/$entry
      -- CP-element group 352: 	 branch_block_stmt_714/whilex_xbody682_ifx_xthen717_PhiReq/$exit
      -- 
    if_choice_transition_6394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2622_branch_ack_1, ack => zeropad3D_CP_2152_elements(352)); -- 
    -- CP-element group 353:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353: 	355 
    -- CP-element group 353: 	357 
    -- CP-element group 353:  members (27) 
      -- CP-element group 353: 	 branch_block_stmt_714/merge_stmt_2628__exit__
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653__entry__
      -- CP-element group 353: 	 branch_block_stmt_714/if_stmt_2622_else_link/$exit
      -- CP-element group 353: 	 branch_block_stmt_714/if_stmt_2622_else_link/else_choice_transition
      -- CP-element group 353: 	 branch_block_stmt_714/whilex_xbody682_lorx_xlhsx_xfalse689
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_update_start_
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_word_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/word_access_start/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/word_access_start/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/word_access_start/word_0/rr
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/word_access_complete/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/word_access_complete/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/word_access_complete/word_0/cr
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_update_start_
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Update/cr
      -- CP-element group 353: 	 branch_block_stmt_714/whilex_xbody682_lorx_xlhsx_xfalse689_PhiReq/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/whilex_xbody682_lorx_xlhsx_xfalse689_PhiReq/$exit
      -- CP-element group 353: 	 branch_block_stmt_714/merge_stmt_2628_PhiReqMerge
      -- CP-element group 353: 	 branch_block_stmt_714/merge_stmt_2628_PhiAck/$entry
      -- CP-element group 353: 	 branch_block_stmt_714/merge_stmt_2628_PhiAck/$exit
      -- CP-element group 353: 	 branch_block_stmt_714/merge_stmt_2628_PhiAck/dummy
      -- 
    else_choice_transition_6398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2622_branch_ack_0, ack => zeropad3D_CP_2152_elements(353)); -- 
    rr_6419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(353), ack => LOAD_row_high_2630_load_0_req_0); -- 
    cr_6430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(353), ack => LOAD_row_high_2630_load_0_req_1); -- 
    cr_6449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(353), ack => type_cast_2634_inst_req_1); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (5) 
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/word_access_start/$exit
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/word_access_start/word_0/$exit
      -- CP-element group 354: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Sample/word_access_start/word_0/ra
      -- 
    ra_6420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2630_load_0_ack_0, ack => zeropad3D_CP_2152_elements(354)); -- 
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (12) 
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/word_access_complete/$exit
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/word_access_complete/word_0/$exit
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/word_access_complete/word_0/ca
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/LOAD_row_high_2630_Merge/$entry
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/LOAD_row_high_2630_Merge/$exit
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/LOAD_row_high_2630_Merge/merge_req
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/LOAD_row_high_2630_Update/LOAD_row_high_2630_Merge/merge_ack
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Sample/rr
      -- 
    ca_6431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2630_load_0_ack_1, ack => zeropad3D_CP_2152_elements(355)); -- 
    rr_6444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(355), ack => type_cast_2634_inst_req_0); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Sample/ra
      -- 
    ra_6445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2634_inst_ack_0, ack => zeropad3D_CP_2152_elements(356)); -- 
    -- CP-element group 357:  branch  transition  place  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	353 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (13) 
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653__exit__
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654__entry__
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/$exit
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_714/assign_stmt_2631_to_assign_stmt_2653/type_cast_2634_Update/ca
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654_dead_link/$entry
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654_eval_test/$entry
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654_eval_test/$exit
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654_eval_test/branch_req
      -- CP-element group 357: 	 branch_block_stmt_714/R_cmp698_2655_place
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654_if_link/$entry
      -- CP-element group 357: 	 branch_block_stmt_714/if_stmt_2654_else_link/$entry
      -- 
    ca_6450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2634_inst_ack_1, ack => zeropad3D_CP_2152_elements(357)); -- 
    branch_req_6458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(357), ack => if_stmt_2654_branch_req_0); -- 
    -- CP-element group 358:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: 	361 
    -- CP-element group 358:  members (18) 
      -- CP-element group 358: 	 branch_block_stmt_714/merge_stmt_2660__exit__
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672__entry__
      -- CP-element group 358: 	 branch_block_stmt_714/if_stmt_2654_if_link/$exit
      -- CP-element group 358: 	 branch_block_stmt_714/if_stmt_2654_if_link/if_choice_transition
      -- CP-element group 358: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_lorx_xlhsx_xfalse700
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/$entry
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_update_start_
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Sample/rr
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Update/$entry
      -- CP-element group 358: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Update/cr
      -- CP-element group 358: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_lorx_xlhsx_xfalse700_PhiReq/$entry
      -- CP-element group 358: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_lorx_xlhsx_xfalse700_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_714/merge_stmt_2660_PhiReqMerge
      -- CP-element group 358: 	 branch_block_stmt_714/merge_stmt_2660_PhiAck/$entry
      -- CP-element group 358: 	 branch_block_stmt_714/merge_stmt_2660_PhiAck/$exit
      -- CP-element group 358: 	 branch_block_stmt_714/merge_stmt_2660_PhiAck/dummy
      -- 
    if_choice_transition_6463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2654_branch_ack_1, ack => zeropad3D_CP_2152_elements(358)); -- 
    rr_6480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(358), ack => type_cast_2664_inst_req_0); -- 
    cr_6485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(358), ack => type_cast_2664_inst_req_1); -- 
    -- CP-element group 359:  transition  place  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	979 
    -- CP-element group 359:  members (5) 
      -- CP-element group 359: 	 branch_block_stmt_714/if_stmt_2654_else_link/$exit
      -- CP-element group 359: 	 branch_block_stmt_714/if_stmt_2654_else_link/else_choice_transition
      -- CP-element group 359: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_ifx_xthen717
      -- CP-element group 359: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_ifx_xthen717_PhiReq/$entry
      -- CP-element group 359: 	 branch_block_stmt_714/lorx_xlhsx_xfalse689_ifx_xthen717_PhiReq/$exit
      -- 
    else_choice_transition_6467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2654_branch_ack_0, ack => zeropad3D_CP_2152_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Sample/ra
      -- 
    ra_6481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2664_inst_ack_0, ack => zeropad3D_CP_2152_elements(360)); -- 
    -- CP-element group 361:  branch  transition  place  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	358 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (13) 
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673__entry__
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672__exit__
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/$exit
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_714/assign_stmt_2665_to_assign_stmt_2672/type_cast_2664_Update/ca
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673_dead_link/$entry
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673_eval_test/$entry
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673_eval_test/$exit
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673_eval_test/branch_req
      -- CP-element group 361: 	 branch_block_stmt_714/R_cmp705_2674_place
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673_if_link/$entry
      -- CP-element group 361: 	 branch_block_stmt_714/if_stmt_2673_else_link/$entry
      -- 
    ca_6486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2664_inst_ack_1, ack => zeropad3D_CP_2152_elements(361)); -- 
    branch_req_6494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(361), ack => if_stmt_2673_branch_req_0); -- 
    -- CP-element group 362:  transition  place  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	979 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 branch_block_stmt_714/if_stmt_2673_if_link/$exit
      -- CP-element group 362: 	 branch_block_stmt_714/if_stmt_2673_if_link/if_choice_transition
      -- CP-element group 362: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_ifx_xthen717
      -- CP-element group 362: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_ifx_xthen717_PhiReq/$entry
      -- CP-element group 362: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_ifx_xthen717_PhiReq/$exit
      -- 
    if_choice_transition_6499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2673_branch_ack_1, ack => zeropad3D_CP_2152_elements(362)); -- 
    -- CP-element group 363:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363: 	365 
    -- CP-element group 363: 	367 
    -- CP-element group 363:  members (27) 
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698__entry__
      -- CP-element group 363: 	 branch_block_stmt_714/merge_stmt_2679__exit__
      -- CP-element group 363: 	 branch_block_stmt_714/if_stmt_2673_else_link/$exit
      -- CP-element group 363: 	 branch_block_stmt_714/if_stmt_2673_else_link/else_choice_transition
      -- CP-element group 363: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_lorx_xlhsx_xfalse707
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_update_start_
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_word_address_calculated
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_root_address_calculated
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/word_access_start/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/word_access_start/word_0/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/word_access_start/word_0/rr
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/word_access_complete/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/word_access_complete/word_0/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/word_access_complete/word_0/cr
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_update_start_
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Update/cr
      -- CP-element group 363: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_lorx_xlhsx_xfalse707_PhiReq/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/lorx_xlhsx_xfalse700_lorx_xlhsx_xfalse707_PhiReq/$exit
      -- CP-element group 363: 	 branch_block_stmt_714/merge_stmt_2679_PhiReqMerge
      -- CP-element group 363: 	 branch_block_stmt_714/merge_stmt_2679_PhiAck/$entry
      -- CP-element group 363: 	 branch_block_stmt_714/merge_stmt_2679_PhiAck/$exit
      -- CP-element group 363: 	 branch_block_stmt_714/merge_stmt_2679_PhiAck/dummy
      -- 
    else_choice_transition_6503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2673_branch_ack_0, ack => zeropad3D_CP_2152_elements(363)); -- 
    rr_6524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(363), ack => LOAD_col_high_2681_load_0_req_0); -- 
    cr_6535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(363), ack => LOAD_col_high_2681_load_0_req_1); -- 
    cr_6554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(363), ack => type_cast_2685_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/word_access_start/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/word_access_start/word_0/$exit
      -- CP-element group 364: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Sample/word_access_start/word_0/ra
      -- 
    ra_6525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2681_load_0_ack_0, ack => zeropad3D_CP_2152_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (12) 
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/word_access_complete/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/word_access_complete/word_0/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/word_access_complete/word_0/ca
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/LOAD_col_high_2681_Merge/$entry
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/LOAD_col_high_2681_Merge/$exit
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/LOAD_col_high_2681_Merge/merge_req
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/LOAD_col_high_2681_Update/LOAD_col_high_2681_Merge/merge_ack
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Sample/rr
      -- 
    ca_6536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2681_load_0_ack_1, ack => zeropad3D_CP_2152_elements(365)); -- 
    rr_6549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(365), ack => type_cast_2685_inst_req_0); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Sample/ra
      -- 
    ra_6550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_0, ack => zeropad3D_CP_2152_elements(366)); -- 
    -- CP-element group 367:  branch  transition  place  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	363 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (13) 
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699__entry__
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698__exit__
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/$exit
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_714/assign_stmt_2682_to_assign_stmt_2698/type_cast_2685_Update/ca
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699_dead_link/$entry
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699_eval_test/$entry
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699_eval_test/$exit
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699_eval_test/branch_req
      -- CP-element group 367: 	 branch_block_stmt_714/R_cmp715_2700_place
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699_if_link/$entry
      -- CP-element group 367: 	 branch_block_stmt_714/if_stmt_2699_else_link/$entry
      -- 
    ca_6555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_1, ack => zeropad3D_CP_2152_elements(367)); -- 
    branch_req_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(367), ack => if_stmt_2699_branch_req_0); -- 
    -- CP-element group 368:  fork  transition  place  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	384 
    -- CP-element group 368: 	385 
    -- CP-element group 368: 	387 
    -- CP-element group 368: 	389 
    -- CP-element group 368: 	391 
    -- CP-element group 368: 	393 
    -- CP-element group 368: 	395 
    -- CP-element group 368: 	397 
    -- CP-element group 368: 	399 
    -- CP-element group 368: 	402 
    -- CP-element group 368:  members (46) 
      -- CP-element group 368: 	 branch_block_stmt_714/merge_stmt_2763__exit__
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868__entry__
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/word_access_complete/word_0/cr
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/word_access_complete/word_0/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_update_start
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_complete/req
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Update/req
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_update_start
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/word_access_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_complete/req
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Sample/rr
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_update_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Update/req
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/if_stmt_2699_if_link/$exit
      -- CP-element group 368: 	 branch_block_stmt_714/if_stmt_2699_if_link/if_choice_transition
      -- CP-element group 368: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xelse738
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/word_access_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/word_access_complete/word_0/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/word_access_complete/word_0/cr
      -- CP-element group 368: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xelse738_PhiReq/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xelse738_PhiReq/$exit
      -- CP-element group 368: 	 branch_block_stmt_714/merge_stmt_2763_PhiReqMerge
      -- CP-element group 368: 	 branch_block_stmt_714/merge_stmt_2763_PhiAck/$entry
      -- CP-element group 368: 	 branch_block_stmt_714/merge_stmt_2763_PhiAck/$exit
      -- CP-element group 368: 	 branch_block_stmt_714/merge_stmt_2763_PhiAck/dummy
      -- 
    if_choice_transition_6568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2699_branch_ack_1, ack => zeropad3D_CP_2152_elements(368)); -- 
    cr_6836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => ptr_deref_2842_load_0_req_1); -- 
    req_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => addr_of_2863_final_reg_req_1); -- 
    cr_6855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => type_cast_2856_inst_req_1); -- 
    req_6776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => array_obj_ref_2837_index_offset_req_1); -- 
    req_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => addr_of_2838_final_reg_req_1); -- 
    cr_6745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => type_cast_2831_inst_req_1); -- 
    cr_6731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => type_cast_2767_inst_req_1); -- 
    rr_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => type_cast_2767_inst_req_0); -- 
    req_6886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => array_obj_ref_2862_index_offset_req_1); -- 
    cr_6951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(368), ack => ptr_deref_2866_store_0_req_1); -- 
    -- CP-element group 369:  transition  place  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	979 
    -- CP-element group 369:  members (5) 
      -- CP-element group 369: 	 branch_block_stmt_714/if_stmt_2699_else_link/$exit
      -- CP-element group 369: 	 branch_block_stmt_714/if_stmt_2699_else_link/else_choice_transition
      -- CP-element group 369: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xthen717
      -- CP-element group 369: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xthen717_PhiReq/$entry
      -- CP-element group 369: 	 branch_block_stmt_714/lorx_xlhsx_xfalse707_ifx_xthen717_PhiReq/$exit
      -- 
    else_choice_transition_6572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2699_branch_ack_0, ack => zeropad3D_CP_2152_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	979 
    -- CP-element group 370: successors 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Sample/ra
      -- 
    ra_6586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => zeropad3D_CP_2152_elements(370)); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	979 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	374 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Update/ca
      -- 
    ca_6591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => zeropad3D_CP_2152_elements(371)); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	979 
    -- CP-element group 372: successors 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Sample/ra
      -- 
    ra_6600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2714_inst_ack_0, ack => zeropad3D_CP_2152_elements(372)); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	979 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Update/ca
      -- 
    ca_6605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2714_inst_ack_1, ack => zeropad3D_CP_2152_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	371 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Sample/rr
      -- 
    rr_6613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(374), ack => type_cast_2748_inst_req_0); -- 
    zeropad3D_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(371) & zeropad3D_CP_2152_elements(373);
      gj_zeropad3D_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Sample/ra
      -- 
    ra_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2748_inst_ack_0, ack => zeropad3D_CP_2152_elements(375)); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	979 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (16) 
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_scale_1/$entry
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_scale_1/$exit
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_scale_1/scale_rename_req
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_scale_1/scale_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_resize_1/index_resize_ack
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_resize_1/index_resize_req
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_resize_1/$exit
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_resize_1/$entry
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Sample/req
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_computed_1
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_scaled_1
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_index_resized_1
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Update/ca
      -- 
    ca_6619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2748_inst_ack_1, ack => zeropad3D_CP_2152_elements(376)); -- 
    req_6644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(376), ack => array_obj_ref_2754_index_offset_req_0); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	383 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_sample_complete
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Sample/ack
      -- CP-element group 377: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Sample/$exit
      -- 
    ack_6645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2754_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(377)); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	979 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (11) 
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_request/$entry
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_request/req
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_base_plus_offset/sum_rename_ack
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_base_plus_offset/sum_rename_req
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_base_plus_offset/$exit
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_base_plus_offset/$entry
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Update/ack
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_root_address_calculated
      -- CP-element group 378: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_offset_calculated
      -- 
    ack_6650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2754_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(378)); -- 
    req_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(378), ack => addr_of_2755_final_reg_req_0); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_request/$exit
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_request/ack
      -- CP-element group 379: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_sample_completed_
      -- 
    ack_6660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2755_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(379)); -- 
    -- CP-element group 380:  join  fork  transition  input  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	979 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (28) 
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_root_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_address_resized
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_addr_resize/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_addr_resize/$exit
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/ptr_deref_2758_Split/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_word_addrgen/root_register_ack
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_word_addrgen/root_register_req
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_word_addrgen/$exit
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_word_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_word_addrgen/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_plus_offset/sum_rename_ack
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_plus_offset/sum_rename_req
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_plus_offset/$exit
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_complete/ack
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_plus_offset/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_addr_resize/base_resize_ack
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/word_access_start/word_0/rr
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_base_addr_resize/base_resize_req
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/word_access_start/word_0/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_complete/$exit
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/word_access_start/$entry
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/ptr_deref_2758_Split/split_ack
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/ptr_deref_2758_Split/split_req
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/ptr_deref_2758_Split/$exit
      -- CP-element group 380: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_update_completed_
      -- 
    ack_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2755_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(380)); -- 
    rr_6703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(380), ack => ptr_deref_2758_store_0_req_0); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/word_access_start/word_0/ra
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/word_access_start/word_0/$exit
      -- CP-element group 381: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Sample/word_access_start/$exit
      -- 
    ra_6704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2758_store_0_ack_0, ack => zeropad3D_CP_2152_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	979 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (5) 
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/word_access_complete/word_0/ca
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/word_access_complete/word_0/$exit
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/word_access_complete/$exit
      -- CP-element group 382: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/$exit
      -- 
    ca_6715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2758_store_0_ack_1, ack => zeropad3D_CP_2152_elements(382)); -- 
    -- CP-element group 383:  join  transition  place  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	377 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	980 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761__exit__
      -- CP-element group 383: 	 branch_block_stmt_714/ifx_xthen717_ifx_xend786
      -- CP-element group 383: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/$exit
      -- CP-element group 383: 	 branch_block_stmt_714/ifx_xthen717_ifx_xend786_PhiReq/$entry
      -- CP-element group 383: 	 branch_block_stmt_714/ifx_xthen717_ifx_xend786_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(377) & zeropad3D_CP_2152_elements(382);
      gj_zeropad3D_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	368 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Sample/ra
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_sample_completed_
      -- 
    ra_6727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_0, ack => zeropad3D_CP_2152_elements(384)); -- 
    -- CP-element group 385:  fork  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	368 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385: 	394 
    -- CP-element group 385:  members (9) 
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Sample/rr
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Sample/rr
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Update/ca
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2767_update_completed_
      -- 
    ca_6732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_1, ack => zeropad3D_CP_2152_elements(385)); -- 
    rr_6740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(385), ack => type_cast_2831_inst_req_0); -- 
    rr_6850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(385), ack => type_cast_2856_inst_req_0); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Sample/ra
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_sample_completed_
      -- 
    ra_6741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2831_inst_ack_0, ack => zeropad3D_CP_2152_elements(386)); -- 
    -- CP-element group 387:  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	368 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (16) 
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Sample/req
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_scale_1/scale_rename_ack
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_scale_1/scale_rename_req
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_scale_1/$exit
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_scale_1/$entry
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_resize_1/index_resize_ack
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_resize_1/index_resize_req
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_resize_1/$exit
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_resize_1/$entry
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_computed_1
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_scaled_1
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_index_resized_1
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Update/ca
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2831_update_completed_
      -- 
    ca_6746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2831_inst_ack_1, ack => zeropad3D_CP_2152_elements(387)); -- 
    req_6771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(387), ack => array_obj_ref_2837_index_offset_req_0); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	403 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Sample/ack
      -- CP-element group 388: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_sample_complete
      -- 
    ack_6772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2837_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(388)); -- 
    -- CP-element group 389:  transition  input  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	368 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (11) 
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_base_plus_offset/$exit
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_base_plus_offset/sum_rename_req
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_base_plus_offset/sum_rename_ack
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_request/$entry
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_request/req
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_base_plus_offset/$entry
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Update/ack
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_final_index_sum_regn_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_offset_calculated
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2837_root_address_calculated
      -- CP-element group 389: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_sample_start_
      -- 
    ack_6777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2837_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(389)); -- 
    req_6786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(389), ack => addr_of_2838_final_reg_req_0); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_request/$exit
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_request/ack
      -- CP-element group 390: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_sample_completed_
      -- 
    ack_6787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2838_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(390)); -- 
    -- CP-element group 391:  join  fork  transition  input  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	368 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (24) 
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_word_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_root_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_address_resized
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_addr_resize/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_complete/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_addr_resize/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/word_access_start/word_0/rr
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_complete/ack
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/word_access_start/word_0/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/word_access_start/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2838_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_word_addrgen/root_register_ack
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_word_addrgen/root_register_req
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_word_addrgen/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_word_addrgen/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_plus_offset/sum_rename_ack
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_plus_offset/sum_rename_req
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_plus_offset/$exit
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_plus_offset/$entry
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_addr_resize/base_resize_ack
      -- CP-element group 391: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_base_addr_resize/base_resize_req
      -- 
    ack_6792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2838_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(391)); -- 
    rr_6825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(391), ack => ptr_deref_2842_load_0_req_0); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (5) 
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/word_access_start/word_0/ra
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/word_access_start/word_0/$exit
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/word_access_start/$exit
      -- CP-element group 392: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Sample/$exit
      -- 
    ra_6826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2842_load_0_ack_0, ack => zeropad3D_CP_2152_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	368 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	400 
    -- CP-element group 393:  members (9) 
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/ptr_deref_2842_Merge/$exit
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/ptr_deref_2842_Merge/merge_req
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/ptr_deref_2842_Merge/merge_ack
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/ptr_deref_2842_Merge/$entry
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/word_access_complete/word_0/ca
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/word_access_complete/word_0/$exit
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/word_access_complete/$exit
      -- CP-element group 393: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2842_Update/$exit
      -- 
    ca_6837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2842_load_0_ack_1, ack => zeropad3D_CP_2152_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	385 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Sample/ra
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_sample_completed_
      -- 
    ra_6851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2856_inst_ack_0, ack => zeropad3D_CP_2152_elements(394)); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	368 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (16) 
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_resized_1
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_scaled_1
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Sample/req
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Update/ca
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_scale_1/scale_rename_ack
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_scale_1/scale_rename_req
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_scale_1/$exit
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_scale_1/$entry
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_resize_1/index_resize_ack
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_resize_1/index_resize_req
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_resize_1/$exit
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_resize_1/$entry
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/type_cast_2856_update_completed_
      -- CP-element group 395: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_index_computed_1
      -- 
    ca_6856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2856_inst_ack_1, ack => zeropad3D_CP_2152_elements(395)); -- 
    req_6881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(395), ack => array_obj_ref_2862_index_offset_req_0); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	403 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Sample/ack
      -- CP-element group 396: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_sample_complete
      -- 
    ack_6882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2862_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(396)); -- 
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	368 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (11) 
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_root_address_calculated
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_offset_calculated
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_request/$entry
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_request/req
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_base_plus_offset/sum_rename_ack
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_base_plus_offset/sum_rename_req
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_base_plus_offset/$exit
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_base_plus_offset/$entry
      -- CP-element group 397: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/array_obj_ref_2862_final_index_sum_regn_Update/ack
      -- 
    ack_6887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2862_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(397)); -- 
    req_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(397), ack => addr_of_2863_final_reg_req_0); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_request/ack
      -- CP-element group 398: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_request/$exit
      -- 
    ack_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2863_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(398)); -- 
    -- CP-element group 399:  fork  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	368 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (19) 
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_address_calculated
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_word_address_calculated
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_root_address_calculated
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_complete/ack
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_address_resized
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_complete/$exit
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_addr_resize/$entry
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_addr_resize/$exit
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/addr_of_2863_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_addr_resize/base_resize_req
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_addr_resize/base_resize_ack
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_plus_offset/$entry
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_plus_offset/$exit
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_plus_offset/sum_rename_req
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_base_plus_offset/sum_rename_ack
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_word_addrgen/$entry
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_word_addrgen/$exit
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_word_addrgen/root_register_req
      -- CP-element group 399: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_word_addrgen/root_register_ack
      -- 
    ack_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2863_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(399)); -- 
    -- CP-element group 400:  join  transition  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	393 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (9) 
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/ptr_deref_2866_Split/$entry
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/ptr_deref_2866_Split/$exit
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/ptr_deref_2866_Split/split_req
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/ptr_deref_2866_Split/split_ack
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/word_access_start/$entry
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/word_access_start/word_0/$entry
      -- CP-element group 400: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/word_access_start/word_0/rr
      -- 
    rr_6940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(400), ack => ptr_deref_2866_store_0_req_0); -- 
    zeropad3D_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(393) & zeropad3D_CP_2152_elements(399);
      gj_zeropad3D_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401:  members (5) 
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_sample_completed_
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/word_access_start/$exit
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/word_access_start/word_0/$exit
      -- CP-element group 401: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Sample/word_access_start/word_0/ra
      -- 
    ra_6941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2866_store_0_ack_0, ack => zeropad3D_CP_2152_elements(401)); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	368 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (5) 
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/word_access_complete/$exit
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/word_access_complete/word_0/$exit
      -- CP-element group 402: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/ptr_deref_2866_Update/word_access_complete/word_0/ca
      -- 
    ca_6952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2866_store_0_ack_1, ack => zeropad3D_CP_2152_elements(402)); -- 
    -- CP-element group 403:  join  transition  place  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	388 
    -- CP-element group 403: 	396 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	980 
    -- CP-element group 403:  members (5) 
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868__exit__
      -- CP-element group 403: 	 branch_block_stmt_714/ifx_xelse738_ifx_xend786
      -- CP-element group 403: 	 branch_block_stmt_714/assign_stmt_2768_to_assign_stmt_2868/$exit
      -- CP-element group 403: 	 branch_block_stmt_714/ifx_xelse738_ifx_xend786_PhiReq/$entry
      -- CP-element group 403: 	 branch_block_stmt_714/ifx_xelse738_ifx_xend786_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_403: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_403"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(388) & zeropad3D_CP_2152_elements(396) & zeropad3D_CP_2152_elements(402);
      gj_zeropad3D_cp_element_group_403 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(403), clk => clk, reset => reset); --
    end block;
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	980 
    -- CP-element group 404: successors 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_sample_completed_
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Sample/ra
      -- 
    ra_6964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2874_inst_ack_0, ack => zeropad3D_CP_2152_elements(404)); -- 
    -- CP-element group 405:  branch  transition  place  input  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	980 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405: 	407 
    -- CP-element group 405:  members (13) 
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889__entry__
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888__exit__
      -- CP-element group 405: 	 branch_block_stmt_714/R_cmp794_2890_place
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/$exit
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_update_completed_
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Update/ca
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889_dead_link/$entry
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889_eval_test/$entry
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889_eval_test/$exit
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889_eval_test/branch_req
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889_if_link/$entry
      -- CP-element group 405: 	 branch_block_stmt_714/if_stmt_2889_else_link/$entry
      -- 
    ca_6969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2874_inst_ack_1, ack => zeropad3D_CP_2152_elements(405)); -- 
    branch_req_6977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(405), ack => if_stmt_2889_branch_req_0); -- 
    -- CP-element group 406:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	989 
    -- CP-element group 406: 	990 
    -- CP-element group 406: 	992 
    -- CP-element group 406: 	993 
    -- CP-element group 406: 	995 
    -- CP-element group 406: 	996 
    -- CP-element group 406:  members (40) 
      -- CP-element group 406: 	 branch_block_stmt_714/merge_stmt_2895__exit__
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2901__entry__
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2901__exit__
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837
      -- CP-element group 406: 	 branch_block_stmt_714/merge_stmt_2895_PhiReqMerge
      -- CP-element group 406: 	 branch_block_stmt_714/merge_stmt_2895_PhiAck/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/merge_stmt_2895_PhiAck/$exit
      -- CP-element group 406: 	 branch_block_stmt_714/merge_stmt_2895_PhiAck/dummy
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xend786_ifx_xthen796
      -- CP-element group 406: 	 branch_block_stmt_714/if_stmt_2889_if_link/$exit
      -- CP-element group 406: 	 branch_block_stmt_714/if_stmt_2889_if_link/if_choice_transition
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2901/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/assign_stmt_2901/$exit
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xend786_ifx_xthen796_PhiReq/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xend786_ifx_xthen796_PhiReq/$exit
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Update/cr
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Update/cr
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2889_branch_ack_1, ack => zeropad3D_CP_2152_elements(406)); -- 
    rr_12890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(406), ack => type_cast_2985_inst_req_0); -- 
    cr_12895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(406), ack => type_cast_2985_inst_req_1); -- 
    rr_12913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(406), ack => type_cast_2992_inst_req_0); -- 
    cr_12918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(406), ack => type_cast_2992_inst_req_1); -- 
    rr_12936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(406), ack => type_cast_2998_inst_req_0); -- 
    cr_12941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(406), ack => type_cast_2998_inst_req_1); -- 
    -- CP-element group 407:  fork  transition  place  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	405 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407: 	409 
    -- CP-element group 407: 	410 
    -- CP-element group 407: 	411 
    -- CP-element group 407: 	413 
    -- CP-element group 407: 	416 
    -- CP-element group 407: 	418 
    -- CP-element group 407: 	419 
    -- CP-element group 407: 	420 
    -- CP-element group 407: 	422 
    -- CP-element group 407:  members (54) 
      -- CP-element group 407: 	 branch_block_stmt_714/merge_stmt_2903__exit__
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974__entry__
      -- CP-element group 407: 	 branch_block_stmt_714/ifx_xend786_ifx_xelse801_PhiReq/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/ifx_xend786_ifx_xelse801_PhiReq/$exit
      -- CP-element group 407: 	 branch_block_stmt_714/ifx_xend786_ifx_xelse801
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2889_else_link/$exit
      -- CP-element group 407: 	 branch_block_stmt_714/if_stmt_2889_else_link/else_choice_transition
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Sample/rr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_word_address_calculated
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_root_address_calculated
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/word_access_start/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/word_access_start/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/word_access_start/word_0/rr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/word_access_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/word_access_complete/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/word_access_complete/word_0/cr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_word_address_calculated
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_root_address_calculated
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/word_access_start/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/word_access_start/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/word_access_start/word_0/rr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/word_access_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/word_access_complete/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/word_access_complete/word_0/cr
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_update_start_
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_714/merge_stmt_2903_PhiReqMerge
      -- CP-element group 407: 	 branch_block_stmt_714/merge_stmt_2903_PhiAck/$entry
      -- CP-element group 407: 	 branch_block_stmt_714/merge_stmt_2903_PhiAck/$exit
      -- CP-element group 407: 	 branch_block_stmt_714/merge_stmt_2903_PhiAck/dummy
      -- 
    else_choice_transition_6986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2889_branch_ack_0, ack => zeropad3D_CP_2152_elements(407)); -- 
    rr_7002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => type_cast_2913_inst_req_0); -- 
    cr_7007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => type_cast_2913_inst_req_1); -- 
    rr_7024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => LOAD_col_high_2916_load_0_req_0); -- 
    cr_7035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => LOAD_col_high_2916_load_0_req_1); -- 
    cr_7054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => type_cast_2920_inst_req_1); -- 
    cr_7068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => type_cast_2934_inst_req_1); -- 
    cr_7082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => type_cast_2950_inst_req_1); -- 
    rr_7099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => LOAD_row_high_2953_load_0_req_0); -- 
    cr_7110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => LOAD_row_high_2953_load_0_req_1); -- 
    cr_7129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(407), ack => type_cast_2957_inst_req_1); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_sample_completed_
      -- CP-element group 408: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Sample/$exit
      -- CP-element group 408: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Sample/ra
      -- 
    ra_7003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_0, ack => zeropad3D_CP_2152_elements(408)); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	407 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	414 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_update_completed_
      -- CP-element group 409: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Update/$exit
      -- CP-element group 409: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2913_Update/ca
      -- 
    ca_7008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2913_inst_ack_1, ack => zeropad3D_CP_2152_elements(409)); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	407 
    -- CP-element group 410: successors 
    -- CP-element group 410:  members (5) 
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/word_access_start/$exit
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/word_access_start/word_0/$exit
      -- CP-element group 410: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Sample/word_access_start/word_0/ra
      -- 
    ra_7025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2916_load_0_ack_0, ack => zeropad3D_CP_2152_elements(410)); -- 
    -- CP-element group 411:  transition  input  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	407 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (12) 
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/word_access_complete/$exit
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/word_access_complete/word_0/$exit
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/word_access_complete/word_0/ca
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/LOAD_col_high_2916_Merge/$entry
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/LOAD_col_high_2916_Merge/$exit
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/LOAD_col_high_2916_Merge/merge_req
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_col_high_2916_Update/LOAD_col_high_2916_Merge/merge_ack
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Sample/rr
      -- 
    ca_7036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_2916_load_0_ack_1, ack => zeropad3D_CP_2152_elements(411)); -- 
    rr_7049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(411), ack => type_cast_2920_inst_req_0); -- 
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Sample/ra
      -- 
    ra_7050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2920_inst_ack_0, ack => zeropad3D_CP_2152_elements(412)); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	407 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2920_Update/ca
      -- 
    ca_7055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2920_inst_ack_1, ack => zeropad3D_CP_2152_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	409 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_sample_start_
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Sample/rr
      -- 
    rr_7063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(414), ack => type_cast_2934_inst_req_0); -- 
    zeropad3D_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(409) & zeropad3D_CP_2152_elements(413);
      gj_zeropad3D_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  transition  input  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_sample_completed_
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Sample/ra
      -- 
    ra_7064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2934_inst_ack_0, ack => zeropad3D_CP_2152_elements(415)); -- 
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	407 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2934_Update/ca
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_sample_start_
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Sample/$entry
      -- CP-element group 416: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Sample/rr
      -- 
    ca_7069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2934_inst_ack_1, ack => zeropad3D_CP_2152_elements(416)); -- 
    rr_7077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(416), ack => type_cast_2950_inst_req_0); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_sample_completed_
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Sample/$exit
      -- CP-element group 417: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Sample/ra
      -- 
    ra_7078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2950_inst_ack_0, ack => zeropad3D_CP_2152_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	407 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	423 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_update_completed_
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Update/$exit
      -- CP-element group 418: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2950_Update/ca
      -- 
    ca_7083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2950_inst_ack_1, ack => zeropad3D_CP_2152_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	407 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_sample_completed_
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/word_access_start/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/word_access_start/word_0/$exit
      -- CP-element group 419: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Sample/word_access_start/word_0/ra
      -- 
    ra_7100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2953_load_0_ack_0, ack => zeropad3D_CP_2152_elements(419)); -- 
    -- CP-element group 420:  transition  input  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	407 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (12) 
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/word_access_complete/$exit
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/word_access_complete/word_0/$exit
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/word_access_complete/word_0/ca
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/LOAD_row_high_2953_Merge/$entry
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/LOAD_row_high_2953_Merge/$exit
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/LOAD_row_high_2953_Merge/merge_req
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/LOAD_row_high_2953_Update/LOAD_row_high_2953_Merge/merge_ack
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_sample_start_
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Sample/rr
      -- 
    ca_7111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_2953_load_0_ack_1, ack => zeropad3D_CP_2152_elements(420)); -- 
    rr_7124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(420), ack => type_cast_2957_inst_req_0); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_sample_completed_
      -- CP-element group 421: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Sample/ra
      -- 
    ra_7125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2957_inst_ack_0, ack => zeropad3D_CP_2152_elements(421)); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	407 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_update_completed_
      -- CP-element group 422: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/type_cast_2957_Update/ca
      -- 
    ca_7130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2957_inst_ack_1, ack => zeropad3D_CP_2152_elements(422)); -- 
    -- CP-element group 423:  branch  join  transition  place  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	418 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423: 	425 
    -- CP-element group 423:  members (10) 
      -- CP-element group 423: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974__exit__
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975__entry__
      -- CP-element group 423: 	 branch_block_stmt_714/assign_stmt_2909_to_assign_stmt_2974/$exit
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975_dead_link/$entry
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975_eval_test/$entry
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975_eval_test/$exit
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975_eval_test/branch_req
      -- CP-element group 423: 	 branch_block_stmt_714/R_cmp828_2976_place
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975_if_link/$entry
      -- CP-element group 423: 	 branch_block_stmt_714/if_stmt_2975_else_link/$entry
      -- 
    branch_req_7138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(423), ack => if_stmt_2975_branch_req_0); -- 
    zeropad3D_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(418) & zeropad3D_CP_2152_elements(422);
      gj_zeropad3D_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	426 
    -- CP-element group 424: 	427 
    -- CP-element group 424: 	429 
    -- CP-element group 424: 	430 
    -- CP-element group 424: 	431 
    -- CP-element group 424: 	432 
    -- CP-element group 424: 	433 
    -- CP-element group 424: 	434 
    -- CP-element group 424: 	435 
    -- CP-element group 424: 	436 
    -- CP-element group 424: 	437 
    -- CP-element group 424: 	438 
    -- CP-element group 424: 	439 
    -- CP-element group 424: 	441 
    -- CP-element group 424: 	443 
    -- CP-element group 424: 	445 
    -- CP-element group 424:  members (124) 
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138__entry__
      -- CP-element group 424: 	 branch_block_stmt_714/merge_stmt_3003__exit__
      -- CP-element group 424: 	 branch_block_stmt_714/if_stmt_2975_if_link/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/if_stmt_2975_if_link/if_choice_transition
      -- CP-element group 424: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_address_resized
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_addr_resize/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_addr_resize/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_addr_resize/base_resize_req
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_addr_resize/base_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_plus_offset/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_plus_offset/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_plus_offset/sum_rename_req
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_base_plus_offset/sum_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_word_addrgen/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_word_addrgen/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_word_addrgen/root_register_req
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_word_addrgen/root_register_ack
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_address_resized
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_addr_resize/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_addr_resize/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_addr_resize/base_resize_req
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_addr_resize/base_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_plus_offset/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_plus_offset/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_plus_offset/sum_rename_req
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_base_plus_offset/sum_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_word_addrgen/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_word_addrgen/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_word_addrgen/root_register_req
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_word_addrgen/root_register_ack
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_update_start_
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/ifx_xelse801_whilex_xend838_PhiReq/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/merge_stmt_3003_PhiReqMerge
      -- CP-element group 424: 	 branch_block_stmt_714/merge_stmt_3003_PhiAck/$entry
      -- CP-element group 424: 	 branch_block_stmt_714/merge_stmt_3003_PhiAck/$exit
      -- CP-element group 424: 	 branch_block_stmt_714/merge_stmt_3003_PhiAck/dummy
      -- 
    if_choice_transition_7143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2975_branch_ack_1, ack => zeropad3D_CP_2152_elements(424)); -- 
    rr_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_row_high_3006_load_0_req_0); -- 
    cr_7179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_row_high_3006_load_0_req_1); -- 
    cr_7198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => type_cast_3010_inst_req_1); -- 
    rr_7215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_pad_3019_load_0_req_0); -- 
    cr_7226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_pad_3019_load_0_req_1); -- 
    rr_7248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_depth_high_3022_load_0_req_0); -- 
    cr_7259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_depth_high_3022_load_0_req_1); -- 
    rr_7281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_col_high_3025_load_0_req_0); -- 
    cr_7292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => LOAD_col_high_3025_load_0_req_1); -- 
    rr_7331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => ptr_deref_3037_load_0_req_0); -- 
    cr_7342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => ptr_deref_3037_load_0_req_1); -- 
    rr_7381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => ptr_deref_3049_load_0_req_0); -- 
    cr_7392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => ptr_deref_3049_load_0_req_1); -- 
    cr_7411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => type_cast_3053_inst_req_1); -- 
    cr_7425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => type_cast_3057_inst_req_1); -- 
    cr_7439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(424), ack => type_cast_3096_inst_req_1); -- 
    -- CP-element group 425:  fork  transition  place  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	423 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	981 
    -- CP-element group 425: 	982 
    -- CP-element group 425: 	983 
    -- CP-element group 425: 	985 
    -- CP-element group 425: 	986 
    -- CP-element group 425:  members (22) 
      -- CP-element group 425: 	 branch_block_stmt_714/if_stmt_2975_else_link/$exit
      -- CP-element group 425: 	 branch_block_stmt_714/if_stmt_2975_else_link/else_choice_transition
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2982/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Sample/rr
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Update/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Update/cr
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Sample/rr
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Update/$entry
      -- CP-element group 425: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2975_branch_ack_0, ack => zeropad3D_CP_2152_elements(425)); -- 
    rr_12841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(425), ack => type_cast_2994_inst_req_0); -- 
    cr_12846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(425), ack => type_cast_2994_inst_req_1); -- 
    rr_12864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_12864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(425), ack => type_cast_3000_inst_req_0); -- 
    cr_12869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_12869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(425), ack => type_cast_3000_inst_req_1); -- 
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	424 
    -- CP-element group 426: successors 
    -- CP-element group 426:  members (5) 
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_sample_completed_
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/word_access_start/$exit
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/word_access_start/word_0/$exit
      -- CP-element group 426: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Sample/word_access_start/word_0/ra
      -- 
    ra_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3006_load_0_ack_0, ack => zeropad3D_CP_2152_elements(426)); -- 
    -- CP-element group 427:  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	424 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (12) 
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/word_access_complete/$exit
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/word_access_complete/word_0/$exit
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/word_access_complete/word_0/ca
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/LOAD_row_high_3006_Merge/$entry
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/LOAD_row_high_3006_Merge/$exit
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/LOAD_row_high_3006_Merge/merge_req
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_row_high_3006_Update/LOAD_row_high_3006_Merge/merge_ack
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Sample/rr
      -- 
    ca_7180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3006_load_0_ack_1, ack => zeropad3D_CP_2152_elements(427)); -- 
    rr_7193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(427), ack => type_cast_3010_inst_req_0); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Sample/ra
      -- 
    ra_7194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3010_inst_ack_0, ack => zeropad3D_CP_2152_elements(428)); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	424 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	446 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3010_Update/ca
      -- 
    ca_7199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3010_inst_ack_1, ack => zeropad3D_CP_2152_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	424 
    -- CP-element group 430: successors 
    -- CP-element group 430:  members (5) 
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_sample_completed_
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/word_access_start/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/word_access_start/word_0/$exit
      -- CP-element group 430: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Sample/word_access_start/word_0/ra
      -- 
    ra_7216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3019_load_0_ack_0, ack => zeropad3D_CP_2152_elements(430)); -- 
    -- CP-element group 431:  transition  input  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	424 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	444 
    -- CP-element group 431:  members (12) 
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_update_completed_
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/word_access_complete/$exit
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/word_access_complete/word_0/$exit
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/word_access_complete/word_0/ca
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/LOAD_pad_3019_Merge/$entry
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/LOAD_pad_3019_Merge/$exit
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/LOAD_pad_3019_Merge/merge_req
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_pad_3019_Update/LOAD_pad_3019_Merge/merge_ack
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_sample_start_
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Sample/$entry
      -- CP-element group 431: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Sample/rr
      -- 
    ca_7227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3019_load_0_ack_1, ack => zeropad3D_CP_2152_elements(431)); -- 
    rr_7434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(431), ack => type_cast_3096_inst_req_0); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	424 
    -- CP-element group 432: successors 
    -- CP-element group 432:  members (5) 
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/word_access_start/$exit
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/word_access_start/word_0/$exit
      -- CP-element group 432: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Sample/word_access_start/word_0/ra
      -- 
    ra_7249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3022_load_0_ack_0, ack => zeropad3D_CP_2152_elements(432)); -- 
    -- CP-element group 433:  transition  input  output  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	424 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	440 
    -- CP-element group 433:  members (12) 
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/word_access_complete/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/word_access_complete/word_0/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/word_access_complete/word_0/ca
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/LOAD_depth_high_3022_Merge/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/LOAD_depth_high_3022_Merge/$exit
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/LOAD_depth_high_3022_Merge/merge_req
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_depth_high_3022_Update/LOAD_depth_high_3022_Merge/merge_ack
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_sample_start_
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Sample/rr
      -- 
    ca_7260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3022_load_0_ack_1, ack => zeropad3D_CP_2152_elements(433)); -- 
    rr_7406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(433), ack => type_cast_3053_inst_req_0); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	424 
    -- CP-element group 434: successors 
    -- CP-element group 434:  members (5) 
      -- CP-element group 434: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_sample_completed_
      -- CP-element group 434: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/word_access_start/$exit
      -- CP-element group 434: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/word_access_start/word_0/$exit
      -- CP-element group 434: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Sample/word_access_start/word_0/ra
      -- 
    ra_7282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3025_load_0_ack_0, ack => zeropad3D_CP_2152_elements(434)); -- 
    -- CP-element group 435:  transition  input  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	424 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	442 
    -- CP-element group 435:  members (12) 
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_update_completed_
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/word_access_complete/$exit
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/word_access_complete/word_0/$exit
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/word_access_complete/word_0/ca
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/LOAD_col_high_3025_Merge/$entry
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/LOAD_col_high_3025_Merge/$exit
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/LOAD_col_high_3025_Merge/merge_req
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/LOAD_col_high_3025_Update/LOAD_col_high_3025_Merge/merge_ack
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_sample_start_
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Sample/$entry
      -- CP-element group 435: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Sample/rr
      -- 
    ca_7293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3025_load_0_ack_1, ack => zeropad3D_CP_2152_elements(435)); -- 
    rr_7420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(435), ack => type_cast_3057_inst_req_0); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	424 
    -- CP-element group 436: successors 
    -- CP-element group 436:  members (5) 
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_sample_completed_
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/word_access_start/$exit
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/word_access_start/word_0/$exit
      -- CP-element group 436: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Sample/word_access_start/word_0/ra
      -- 
    ra_7332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3037_load_0_ack_0, ack => zeropad3D_CP_2152_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	424 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	446 
    -- CP-element group 437:  members (9) 
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/$exit
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/word_access_complete/$exit
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/word_access_complete/word_0/$exit
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/word_access_complete/word_0/ca
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/ptr_deref_3037_Merge/$entry
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/ptr_deref_3037_Merge/$exit
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/ptr_deref_3037_Merge/merge_req
      -- CP-element group 437: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3037_Update/ptr_deref_3037_Merge/merge_ack
      -- 
    ca_7343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3037_load_0_ack_1, ack => zeropad3D_CP_2152_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	424 
    -- CP-element group 438: successors 
    -- CP-element group 438:  members (5) 
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_sample_completed_
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/word_access_start/$exit
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/word_access_start/word_0/$exit
      -- CP-element group 438: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Sample/word_access_start/word_0/ra
      -- 
    ra_7382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3049_load_0_ack_0, ack => zeropad3D_CP_2152_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	424 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	446 
    -- CP-element group 439:  members (9) 
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_update_completed_
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/word_access_complete/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/word_access_complete/word_0/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/word_access_complete/word_0/ca
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/ptr_deref_3049_Merge/$entry
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/ptr_deref_3049_Merge/$exit
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/ptr_deref_3049_Merge/merge_req
      -- CP-element group 439: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/ptr_deref_3049_Update/ptr_deref_3049_Merge/merge_ack
      -- 
    ca_7393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3049_load_0_ack_1, ack => zeropad3D_CP_2152_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	433 
    -- CP-element group 440: successors 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_sample_completed_
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Sample/ra
      -- 
    ra_7407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3053_inst_ack_0, ack => zeropad3D_CP_2152_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	424 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	446 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_update_completed_
      -- CP-element group 441: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3053_Update/ca
      -- 
    ca_7412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3053_inst_ack_1, ack => zeropad3D_CP_2152_elements(441)); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	435 
    -- CP-element group 442: successors 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_sample_completed_
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Sample/$exit
      -- CP-element group 442: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Sample/ra
      -- 
    ra_7421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3057_inst_ack_0, ack => zeropad3D_CP_2152_elements(442)); -- 
    -- CP-element group 443:  transition  input  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	424 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	446 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_update_completed_
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Update/$exit
      -- CP-element group 443: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3057_Update/ca
      -- 
    ca_7426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3057_inst_ack_1, ack => zeropad3D_CP_2152_elements(443)); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	431 
    -- CP-element group 444: successors 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_sample_completed_
      -- CP-element group 444: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Sample/ra
      -- 
    ra_7435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3096_inst_ack_0, ack => zeropad3D_CP_2152_elements(444)); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	424 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_update_completed_
      -- CP-element group 445: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/type_cast_3096_Update/ca
      -- 
    ca_7440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3096_inst_ack_1, ack => zeropad3D_CP_2152_elements(445)); -- 
    -- CP-element group 446:  join  fork  transition  place  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	429 
    -- CP-element group 446: 	437 
    -- CP-element group 446: 	439 
    -- CP-element group 446: 	441 
    -- CP-element group 446: 	443 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	1014 
    -- CP-element group 446: 	1015 
    -- CP-element group 446: 	1016 
    -- CP-element group 446: 	1018 
    -- CP-element group 446:  members (16) 
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898
      -- CP-element group 446: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138__exit__
      -- CP-element group 446: 	 branch_block_stmt_714/assign_stmt_3007_to_assign_stmt_3138/$exit
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3154/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Sample/rr
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Update/cr
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3141/$entry
      -- CP-element group 446: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/$entry
      -- 
    rr_13057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(446), ack => type_cast_3151_inst_req_0); -- 
    cr_13062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(446), ack => type_cast_3151_inst_req_1); -- 
    zeropad3D_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(429) & zeropad3D_CP_2152_elements(437) & zeropad3D_CP_2152_elements(439) & zeropad3D_CP_2152_elements(441) & zeropad3D_CP_2152_elements(443) & zeropad3D_CP_2152_elements(445);
      gj_zeropad3D_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	1024 
    -- CP-element group 447: successors 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Sample/ra
      -- 
    ra_7452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3165_inst_ack_0, ack => zeropad3D_CP_2152_elements(447)); -- 
    -- CP-element group 448:  branch  transition  place  input  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	1024 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448: 	450 
    -- CP-element group 448:  members (13) 
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174__entry__
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173__exit__
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/$exit
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Update/ca
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174_dead_link/$entry
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174_eval_test/$entry
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174_eval_test/$exit
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174_eval_test/branch_req
      -- CP-element group 448: 	 branch_block_stmt_714/R_cmp903_3175_place
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174_if_link/$entry
      -- CP-element group 448: 	 branch_block_stmt_714/if_stmt_3174_else_link/$entry
      -- 
    ca_7457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3165_inst_ack_1, ack => zeropad3D_CP_2152_elements(448)); -- 
    branch_req_7465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(448), ack => if_stmt_3174_branch_req_0); -- 
    -- CP-element group 449:  transition  place  input  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	1025 
    -- CP-element group 449:  members (5) 
      -- CP-element group 449: 	 branch_block_stmt_714/if_stmt_3174_if_link/$exit
      -- CP-element group 449: 	 branch_block_stmt_714/if_stmt_3174_if_link/if_choice_transition
      -- CP-element group 449: 	 branch_block_stmt_714/whilex_xbody898_ifx_xthen935
      -- CP-element group 449: 	 branch_block_stmt_714/whilex_xbody898_ifx_xthen935_PhiReq/$entry
      -- CP-element group 449: 	 branch_block_stmt_714/whilex_xbody898_ifx_xthen935_PhiReq/$exit
      -- 
    if_choice_transition_7470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3174_branch_ack_1, ack => zeropad3D_CP_2152_elements(449)); -- 
    -- CP-element group 450:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	448 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450: 	452 
    -- CP-element group 450: 	454 
    -- CP-element group 450:  members (27) 
      -- CP-element group 450: 	 branch_block_stmt_714/merge_stmt_3180__exit__
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211__entry__
      -- CP-element group 450: 	 branch_block_stmt_714/if_stmt_3174_else_link/$exit
      -- CP-element group 450: 	 branch_block_stmt_714/if_stmt_3174_else_link/else_choice_transition
      -- CP-element group 450: 	 branch_block_stmt_714/whilex_xbody898_lorx_xlhsx_xfalse905
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_sample_start_
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_update_start_
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_word_address_calculated
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_root_address_calculated
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/word_access_start/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/word_access_start/word_0/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/word_access_start/word_0/rr
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/word_access_complete/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/word_access_complete/word_0/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/word_access_complete/word_0/cr
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_update_start_
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Update/cr
      -- CP-element group 450: 	 branch_block_stmt_714/whilex_xbody898_lorx_xlhsx_xfalse905_PhiReq/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/whilex_xbody898_lorx_xlhsx_xfalse905_PhiReq/$exit
      -- CP-element group 450: 	 branch_block_stmt_714/merge_stmt_3180_PhiReqMerge
      -- CP-element group 450: 	 branch_block_stmt_714/merge_stmt_3180_PhiAck/$entry
      -- CP-element group 450: 	 branch_block_stmt_714/merge_stmt_3180_PhiAck/$exit
      -- CP-element group 450: 	 branch_block_stmt_714/merge_stmt_3180_PhiAck/dummy
      -- 
    else_choice_transition_7474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3174_branch_ack_0, ack => zeropad3D_CP_2152_elements(450)); -- 
    rr_7495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(450), ack => LOAD_row_high_3182_load_0_req_0); -- 
    cr_7506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(450), ack => LOAD_row_high_3182_load_0_req_1); -- 
    cr_7525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(450), ack => type_cast_3186_inst_req_1); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451:  members (5) 
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_sample_completed_
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/word_access_start/$exit
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/word_access_start/word_0/$exit
      -- CP-element group 451: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Sample/word_access_start/word_0/ra
      -- 
    ra_7496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3182_load_0_ack_0, ack => zeropad3D_CP_2152_elements(451)); -- 
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (12) 
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_update_completed_
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/word_access_complete/$exit
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/word_access_complete/word_0/$exit
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/word_access_complete/word_0/ca
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/LOAD_row_high_3182_Merge/$entry
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/LOAD_row_high_3182_Merge/$exit
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/LOAD_row_high_3182_Merge/merge_req
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/LOAD_row_high_3182_Update/LOAD_row_high_3182_Merge/merge_ack
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Sample/rr
      -- 
    ca_7507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3182_load_0_ack_1, ack => zeropad3D_CP_2152_elements(452)); -- 
    rr_7520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(452), ack => type_cast_3186_inst_req_0); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_sample_completed_
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Sample/$exit
      -- CP-element group 453: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Sample/ra
      -- 
    ra_7521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3186_inst_ack_0, ack => zeropad3D_CP_2152_elements(453)); -- 
    -- CP-element group 454:  branch  transition  place  input  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	450 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (13) 
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211__exit__
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212__entry__
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/$exit
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_update_completed_
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Update/$exit
      -- CP-element group 454: 	 branch_block_stmt_714/assign_stmt_3183_to_assign_stmt_3211/type_cast_3186_Update/ca
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212_dead_link/$entry
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212_eval_test/$entry
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212_eval_test/$exit
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212_eval_test/branch_req
      -- CP-element group 454: 	 branch_block_stmt_714/R_cmp915_3213_place
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212_if_link/$entry
      -- CP-element group 454: 	 branch_block_stmt_714/if_stmt_3212_else_link/$entry
      -- 
    ca_7526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3186_inst_ack_1, ack => zeropad3D_CP_2152_elements(454)); -- 
    branch_req_7534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(454), ack => if_stmt_3212_branch_req_0); -- 
    -- CP-element group 455:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	457 
    -- CP-element group 455: 	458 
    -- CP-element group 455:  members (18) 
      -- CP-element group 455: 	 branch_block_stmt_714/merge_stmt_3218__exit__
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230__entry__
      -- CP-element group 455: 	 branch_block_stmt_714/if_stmt_3212_if_link/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/if_stmt_3212_if_link/if_choice_transition
      -- CP-element group 455: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_lorx_xlhsx_xfalse917
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_sample_start_
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_update_start_
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Sample/rr
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_lorx_xlhsx_xfalse917_PhiReq/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_lorx_xlhsx_xfalse917_PhiReq/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/merge_stmt_3218_PhiReqMerge
      -- CP-element group 455: 	 branch_block_stmt_714/merge_stmt_3218_PhiAck/$entry
      -- CP-element group 455: 	 branch_block_stmt_714/merge_stmt_3218_PhiAck/$exit
      -- CP-element group 455: 	 branch_block_stmt_714/merge_stmt_3218_PhiAck/dummy
      -- 
    if_choice_transition_7539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3212_branch_ack_1, ack => zeropad3D_CP_2152_elements(455)); -- 
    rr_7556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(455), ack => type_cast_3222_inst_req_0); -- 
    cr_7561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(455), ack => type_cast_3222_inst_req_1); -- 
    -- CP-element group 456:  transition  place  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	1025 
    -- CP-element group 456:  members (5) 
      -- CP-element group 456: 	 branch_block_stmt_714/if_stmt_3212_else_link/$exit
      -- CP-element group 456: 	 branch_block_stmt_714/if_stmt_3212_else_link/else_choice_transition
      -- CP-element group 456: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_ifx_xthen935
      -- CP-element group 456: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_ifx_xthen935_PhiReq/$entry
      -- CP-element group 456: 	 branch_block_stmt_714/lorx_xlhsx_xfalse905_ifx_xthen935_PhiReq/$exit
      -- 
    else_choice_transition_7543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3212_branch_ack_0, ack => zeropad3D_CP_2152_elements(456)); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	455 
    -- CP-element group 457: successors 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_sample_completed_
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Sample/$exit
      -- CP-element group 457: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Sample/ra
      -- 
    ra_7557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3222_inst_ack_0, ack => zeropad3D_CP_2152_elements(457)); -- 
    -- CP-element group 458:  branch  transition  place  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	455 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458: 	460 
    -- CP-element group 458:  members (13) 
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230__exit__
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231__entry__
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/$exit
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_update_completed_
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Update/$exit
      -- CP-element group 458: 	 branch_block_stmt_714/assign_stmt_3223_to_assign_stmt_3230/type_cast_3222_Update/ca
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231_dead_link/$entry
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231_eval_test/$entry
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231_eval_test/$exit
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231_eval_test/branch_req
      -- CP-element group 458: 	 branch_block_stmt_714/R_cmp922_3232_place
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231_if_link/$entry
      -- CP-element group 458: 	 branch_block_stmt_714/if_stmt_3231_else_link/$entry
      -- 
    ca_7562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3222_inst_ack_1, ack => zeropad3D_CP_2152_elements(458)); -- 
    branch_req_7570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(458), ack => if_stmt_3231_branch_req_0); -- 
    -- CP-element group 459:  transition  place  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	1025 
    -- CP-element group 459:  members (5) 
      -- CP-element group 459: 	 branch_block_stmt_714/if_stmt_3231_if_link/$exit
      -- CP-element group 459: 	 branch_block_stmt_714/if_stmt_3231_if_link/if_choice_transition
      -- CP-element group 459: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_ifx_xthen935
      -- CP-element group 459: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_ifx_xthen935_PhiReq/$entry
      -- CP-element group 459: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_ifx_xthen935_PhiReq/$exit
      -- 
    if_choice_transition_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3231_branch_ack_1, ack => zeropad3D_CP_2152_elements(459)); -- 
    -- CP-element group 460:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460: 	462 
    -- CP-element group 460: 	464 
    -- CP-element group 460:  members (27) 
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262__entry__
      -- CP-element group 460: 	 branch_block_stmt_714/merge_stmt_3237__exit__
      -- CP-element group 460: 	 branch_block_stmt_714/if_stmt_3231_else_link/$exit
      -- CP-element group 460: 	 branch_block_stmt_714/if_stmt_3231_else_link/else_choice_transition
      -- CP-element group 460: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_lorx_xlhsx_xfalse924
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_update_start_
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_word_address_calculated
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_root_address_calculated
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/word_access_start/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/word_access_start/word_0/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/word_access_start/word_0/rr
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/word_access_complete/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/word_access_complete/word_0/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/word_access_complete/word_0/cr
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_update_start_
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Update/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Update/cr
      -- CP-element group 460: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_lorx_xlhsx_xfalse924_PhiReq/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/lorx_xlhsx_xfalse917_lorx_xlhsx_xfalse924_PhiReq/$exit
      -- CP-element group 460: 	 branch_block_stmt_714/merge_stmt_3237_PhiReqMerge
      -- CP-element group 460: 	 branch_block_stmt_714/merge_stmt_3237_PhiAck/$entry
      -- CP-element group 460: 	 branch_block_stmt_714/merge_stmt_3237_PhiAck/$exit
      -- CP-element group 460: 	 branch_block_stmt_714/merge_stmt_3237_PhiAck/dummy
      -- 
    else_choice_transition_7579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3231_branch_ack_0, ack => zeropad3D_CP_2152_elements(460)); -- 
    rr_7600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(460), ack => LOAD_col_high_3239_load_0_req_0); -- 
    cr_7611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(460), ack => LOAD_col_high_3239_load_0_req_1); -- 
    cr_7630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(460), ack => type_cast_3243_inst_req_1); -- 
    -- CP-element group 461:  transition  input  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461:  members (5) 
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/word_access_start/$exit
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/word_access_start/word_0/$exit
      -- CP-element group 461: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Sample/word_access_start/word_0/ra
      -- 
    ra_7601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3239_load_0_ack_0, ack => zeropad3D_CP_2152_elements(461)); -- 
    -- CP-element group 462:  transition  input  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	460 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (12) 
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/word_access_complete/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/word_access_complete/word_0/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/word_access_complete/word_0/ca
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/LOAD_col_high_3239_Merge/$entry
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/LOAD_col_high_3239_Merge/$exit
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/LOAD_col_high_3239_Merge/merge_req
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/LOAD_col_high_3239_Update/LOAD_col_high_3239_Merge/merge_ack
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_sample_start_
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Sample/rr
      -- 
    ca_7612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3239_load_0_ack_1, ack => zeropad3D_CP_2152_elements(462)); -- 
    rr_7625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(462), ack => type_cast_3243_inst_req_0); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_sample_completed_
      -- CP-element group 463: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Sample/ra
      -- 
    ra_7626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3243_inst_ack_0, ack => zeropad3D_CP_2152_elements(463)); -- 
    -- CP-element group 464:  branch  transition  place  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	460 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464: 	466 
    -- CP-element group 464:  members (13) 
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263__entry__
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262__exit__
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/$exit
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_update_completed_
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Update/$exit
      -- CP-element group 464: 	 branch_block_stmt_714/assign_stmt_3240_to_assign_stmt_3262/type_cast_3243_Update/ca
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263_dead_link/$entry
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263_eval_test/$entry
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263_eval_test/$exit
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263_eval_test/branch_req
      -- CP-element group 464: 	 branch_block_stmt_714/R_cmp933_3264_place
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263_if_link/$entry
      -- CP-element group 464: 	 branch_block_stmt_714/if_stmt_3263_else_link/$entry
      -- 
    ca_7631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3243_inst_ack_1, ack => zeropad3D_CP_2152_elements(464)); -- 
    branch_req_7639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(464), ack => if_stmt_3263_branch_req_0); -- 
    -- CP-element group 465:  fork  transition  place  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	481 
    -- CP-element group 465: 	482 
    -- CP-element group 465: 	484 
    -- CP-element group 465: 	486 
    -- CP-element group 465: 	488 
    -- CP-element group 465: 	490 
    -- CP-element group 465: 	492 
    -- CP-element group 465: 	494 
    -- CP-element group 465: 	496 
    -- CP-element group 465: 	499 
    -- CP-element group 465:  members (46) 
      -- CP-element group 465: 	 branch_block_stmt_714/merge_stmt_3327__exit__
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432__entry__
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Update/req
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/word_access_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/word_access_complete/word_0/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/word_access_complete/word_0/cr
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_complete/req
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_update_start
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_complete/req
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Update/req
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_update_start
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_update_start_
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/if_stmt_3263_if_link/$exit
      -- CP-element group 465: 	 branch_block_stmt_714/if_stmt_3263_if_link/if_choice_transition
      -- CP-element group 465: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xelse956
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/word_access_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/word_access_complete/word_0/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/word_access_complete/word_0/cr
      -- CP-element group 465: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xelse956_PhiReq/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xelse956_PhiReq/$exit
      -- CP-element group 465: 	 branch_block_stmt_714/merge_stmt_3327_PhiReqMerge
      -- CP-element group 465: 	 branch_block_stmt_714/merge_stmt_3327_PhiAck/$entry
      -- CP-element group 465: 	 branch_block_stmt_714/merge_stmt_3327_PhiAck/$exit
      -- CP-element group 465: 	 branch_block_stmt_714/merge_stmt_3327_PhiAck/dummy
      -- 
    if_choice_transition_7644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3263_branch_ack_1, ack => zeropad3D_CP_2152_elements(465)); -- 
    req_7962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => array_obj_ref_3426_index_offset_req_1); -- 
    cr_7912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => ptr_deref_3406_load_0_req_1); -- 
    cr_7807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => type_cast_3331_inst_req_1); -- 
    cr_7931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => type_cast_3420_inst_req_1); -- 
    req_7977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => addr_of_3427_final_reg_req_1); -- 
    cr_7821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => type_cast_3395_inst_req_1); -- 
    rr_7802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => type_cast_3331_inst_req_0); -- 
    req_7867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => addr_of_3402_final_reg_req_1); -- 
    req_7852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => array_obj_ref_3401_index_offset_req_1); -- 
    cr_8027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(465), ack => ptr_deref_3430_store_0_req_1); -- 
    -- CP-element group 466:  transition  place  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	464 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	1025 
    -- CP-element group 466:  members (5) 
      -- CP-element group 466: 	 branch_block_stmt_714/if_stmt_3263_else_link/$exit
      -- CP-element group 466: 	 branch_block_stmt_714/if_stmt_3263_else_link/else_choice_transition
      -- CP-element group 466: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xthen935
      -- CP-element group 466: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xthen935_PhiReq/$entry
      -- CP-element group 466: 	 branch_block_stmt_714/lorx_xlhsx_xfalse924_ifx_xthen935_PhiReq/$exit
      -- 
    else_choice_transition_7648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3263_branch_ack_0, ack => zeropad3D_CP_2152_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	1025 
    -- CP-element group 467: successors 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_sample_completed_
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Sample/ra
      -- 
    ra_7662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3273_inst_ack_0, ack => zeropad3D_CP_2152_elements(467)); -- 
    -- CP-element group 468:  transition  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	1025 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	471 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Update/ca
      -- 
    ca_7667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3273_inst_ack_1, ack => zeropad3D_CP_2152_elements(468)); -- 
    -- CP-element group 469:  transition  input  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	1025 
    -- CP-element group 469: successors 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_sample_completed_
      -- CP-element group 469: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Sample/$exit
      -- CP-element group 469: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Sample/ra
      -- 
    ra_7676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3278_inst_ack_0, ack => zeropad3D_CP_2152_elements(469)); -- 
    -- CP-element group 470:  transition  input  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	1025 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_update_completed_
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Update/$exit
      -- CP-element group 470: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Update/ca
      -- 
    ca_7681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3278_inst_ack_1, ack => zeropad3D_CP_2152_elements(470)); -- 
    -- CP-element group 471:  join  transition  output  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	468 
    -- CP-element group 471: 	470 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	472 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_sample_start_
      -- CP-element group 471: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Sample/$entry
      -- CP-element group 471: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Sample/rr
      -- 
    rr_7689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(471), ack => type_cast_3312_inst_req_0); -- 
    zeropad3D_cp_element_group_471: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_471"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(468) & zeropad3D_CP_2152_elements(470);
      gj_zeropad3D_cp_element_group_471 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	471 
    -- CP-element group 472: successors 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_sample_completed_
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Sample/ra
      -- 
    ra_7690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3312_inst_ack_0, ack => zeropad3D_CP_2152_elements(472)); -- 
    -- CP-element group 473:  transition  input  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	1025 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (16) 
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_update_completed_
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Update/ca
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_resized_1
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_scaled_1
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_computed_1
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_resize_1/$entry
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_resize_1/$exit
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_resize_1/index_resize_req
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_resize_1/index_resize_ack
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_scale_1/$entry
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_scale_1/$exit
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_scale_1/scale_rename_req
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_index_scale_1/scale_rename_ack
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Sample/$entry
      -- CP-element group 473: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Sample/req
      -- 
    ca_7695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3312_inst_ack_1, ack => zeropad3D_CP_2152_elements(473)); -- 
    req_7720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(473), ack => array_obj_ref_3318_index_offset_req_0); -- 
    -- CP-element group 474:  transition  input  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	480 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_sample_complete
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Sample/$exit
      -- CP-element group 474: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Sample/ack
      -- 
    ack_7721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3318_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(474)); -- 
    -- CP-element group 475:  transition  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	1025 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (11) 
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_root_address_calculated
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_offset_calculated
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Update/$exit
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Update/ack
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_base_plus_offset/$entry
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_base_plus_offset/$exit
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_base_plus_offset/sum_rename_req
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_base_plus_offset/sum_rename_ack
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_request/$entry
      -- CP-element group 475: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_request/req
      -- 
    ack_7726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3318_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(475)); -- 
    req_7735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(475), ack => addr_of_3319_final_reg_req_0); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_sample_completed_
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_request/$exit
      -- CP-element group 476: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_request/ack
      -- 
    ack_7736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3319_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(476)); -- 
    -- CP-element group 477:  join  fork  transition  input  output  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	1025 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	478 
    -- CP-element group 477:  members (28) 
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/word_access_start/word_0/rr
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/word_access_start/word_0/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/word_access_start/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/ptr_deref_3322_Split/split_ack
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/ptr_deref_3322_Split/split_req
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_update_completed_
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_complete/$exit
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_complete/ack
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_sample_start_
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_address_calculated
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_word_address_calculated
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_root_address_calculated
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_address_resized
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_addr_resize/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_addr_resize/$exit
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_addr_resize/base_resize_req
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_addr_resize/base_resize_ack
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_plus_offset/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_plus_offset/$exit
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_plus_offset/sum_rename_req
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_base_plus_offset/sum_rename_ack
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_word_addrgen/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_word_addrgen/$exit
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_word_addrgen/root_register_req
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_word_addrgen/root_register_ack
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/ptr_deref_3322_Split/$entry
      -- CP-element group 477: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/ptr_deref_3322_Split/$exit
      -- 
    ack_7741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3319_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(477)); -- 
    rr_7779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(477), ack => ptr_deref_3322_store_0_req_0); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	477 
    -- CP-element group 478: successors 
    -- CP-element group 478:  members (5) 
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/word_access_start/word_0/$exit
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/word_access_start/word_0/ra
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/word_access_start/$exit
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_sample_completed_
      -- CP-element group 478: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Sample/$exit
      -- 
    ra_7780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3322_store_0_ack_0, ack => zeropad3D_CP_2152_elements(478)); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	1025 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (5) 
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/word_access_complete/$exit
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/word_access_complete/word_0/$exit
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/word_access_complete/word_0/ca
      -- CP-element group 479: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_update_completed_
      -- 
    ca_7791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3322_store_0_ack_1, ack => zeropad3D_CP_2152_elements(479)); -- 
    -- CP-element group 480:  join  transition  place  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	474 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	1026 
    -- CP-element group 480:  members (5) 
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325__exit__
      -- CP-element group 480: 	 branch_block_stmt_714/ifx_xthen935_ifx_xend1004
      -- CP-element group 480: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/$exit
      -- CP-element group 480: 	 branch_block_stmt_714/ifx_xthen935_ifx_xend1004_PhiReq/$entry
      -- CP-element group 480: 	 branch_block_stmt_714/ifx_xthen935_ifx_xend1004_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_480"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(474) & zeropad3D_CP_2152_elements(479);
      gj_zeropad3D_cp_element_group_480 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481:  transition  input  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	465 
    -- CP-element group 481: successors 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Sample/ra
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Sample/$exit
      -- CP-element group 481: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_sample_completed_
      -- 
    ra_7803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3331_inst_ack_0, ack => zeropad3D_CP_2152_elements(481)); -- 
    -- CP-element group 482:  fork  transition  input  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	465 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482: 	491 
    -- CP-element group 482:  members (9) 
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Update/$exit
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_Update/ca
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3331_update_completed_
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Sample/$entry
      -- 
    ca_7808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3331_inst_ack_1, ack => zeropad3D_CP_2152_elements(482)); -- 
    rr_7816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3395_inst_req_0); -- 
    rr_7926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(482), ack => type_cast_3420_inst_req_0); -- 
    -- CP-element group 483:  transition  input  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Sample/ra
      -- CP-element group 483: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_sample_completed_
      -- 
    ra_7817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3395_inst_ack_0, ack => zeropad3D_CP_2152_elements(483)); -- 
    -- CP-element group 484:  transition  input  output  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	465 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	485 
    -- CP-element group 484:  members (16) 
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Update/ca
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_resize_1/$exit
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_resize_1/index_resize_req
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_resize_1/index_resize_ack
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_scale_1/$entry
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_scale_1/$exit
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_scale_1/scale_rename_req
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_resize_1/$entry
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_computed_1
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_scaled_1
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_resized_1
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Sample/req
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3395_update_completed_
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Sample/$entry
      -- CP-element group 484: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_index_scale_1/scale_rename_ack
      -- 
    ca_7822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3395_inst_ack_1, ack => zeropad3D_CP_2152_elements(484)); -- 
    req_7847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(484), ack => array_obj_ref_3401_index_offset_req_0); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	484 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	500 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Sample/ack
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_sample_complete
      -- 
    ack_7848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3401_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(485)); -- 
    -- CP-element group 486:  transition  input  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	465 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (11) 
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_request/req
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_offset_calculated
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_request/$entry
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_base_plus_offset/sum_rename_ack
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_root_address_calculated
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_base_plus_offset/sum_rename_req
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_base_plus_offset/$exit
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_base_plus_offset/$entry
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Update/ack
      -- CP-element group 486: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3401_final_index_sum_regn_Update/$exit
      -- 
    ack_7853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3401_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(486)); -- 
    req_7862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(486), ack => addr_of_3402_final_reg_req_0); -- 
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_request/ack
      -- CP-element group 487: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_request/$exit
      -- 
    ack_7863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3402_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(487)); -- 
    -- CP-element group 488:  join  fork  transition  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	465 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (24) 
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/word_access_start/word_0/rr
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/word_access_start/word_0/$entry
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/word_access_start/$entry
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_word_addrgen/root_register_ack
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_word_addrgen/root_register_req
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_word_addrgen/$exit
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_word_addrgen/$entry
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_plus_offset/sum_rename_ack
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_plus_offset/sum_rename_req
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_plus_offset/$exit
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_plus_offset/$entry
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_addr_resize/base_resize_ack
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_addr_resize/base_resize_req
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_addr_resize/$exit
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_addr_resize/$entry
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_address_resized
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_root_address_calculated
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_word_address_calculated
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_base_address_calculated
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_sample_start_
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_complete/ack
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_complete/$exit
      -- CP-element group 488: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3402_update_completed_
      -- 
    ack_7868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3402_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(488)); -- 
    rr_7901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(488), ack => ptr_deref_3406_load_0_req_0); -- 
    -- CP-element group 489:  transition  input  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489:  members (5) 
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/word_access_start/word_0/ra
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/word_access_start/word_0/$exit
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/word_access_start/$exit
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_sample_completed_
      -- 
    ra_7902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3406_load_0_ack_0, ack => zeropad3D_CP_2152_elements(489)); -- 
    -- CP-element group 490:  transition  input  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	465 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	497 
    -- CP-element group 490:  members (9) 
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/word_access_complete/$exit
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/word_access_complete/word_0/$exit
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/word_access_complete/word_0/ca
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/ptr_deref_3406_Merge/$entry
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/ptr_deref_3406_Merge/$exit
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/ptr_deref_3406_Merge/merge_req
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/ptr_deref_3406_Merge/merge_ack
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3406_update_completed_
      -- 
    ca_7913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3406_load_0_ack_1, ack => zeropad3D_CP_2152_elements(490)); -- 
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	482 
    -- CP-element group 491: successors 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Sample/ra
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Sample/$exit
      -- 
    ra_7927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3420_inst_ack_0, ack => zeropad3D_CP_2152_elements(491)); -- 
    -- CP-element group 492:  transition  input  output  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	465 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (16) 
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Sample/req
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_scale_1/$exit
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_scale_1/scale_rename_req
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_scale_1/$entry
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_resize_1/index_resize_ack
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_resize_1/index_resize_req
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_resize_1/$exit
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_resize_1/$entry
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_computed_1
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_scaled_1
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_resized_1
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Sample/$entry
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_index_scale_1/scale_rename_ack
      -- CP-element group 492: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/type_cast_3420_Update/ca
      -- 
    ca_7932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3420_inst_ack_1, ack => zeropad3D_CP_2152_elements(492)); -- 
    req_7957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(492), ack => array_obj_ref_3426_index_offset_req_0); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	500 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Sample/ack
      -- CP-element group 493: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Sample/$exit
      -- CP-element group 493: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_sample_complete
      -- 
    ack_7958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3426_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(493)); -- 
    -- CP-element group 494:  transition  input  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	465 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (11) 
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Update/ack
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_base_plus_offset/$entry
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_base_plus_offset/$exit
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_final_index_sum_regn_Update/$exit
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_base_plus_offset/sum_rename_req
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_request/$entry
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_request/req
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_offset_calculated
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_root_address_calculated
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/array_obj_ref_3426_base_plus_offset/sum_rename_ack
      -- CP-element group 494: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_sample_start_
      -- 
    ack_7963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3426_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(494)); -- 
    req_7972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(494), ack => addr_of_3427_final_reg_req_0); -- 
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_request/ack
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_request/$exit
      -- CP-element group 495: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_sample_completed_
      -- 
    ack_7973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3427_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(495)); -- 
    -- CP-element group 496:  fork  transition  input  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	465 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (19) 
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_complete/ack
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_address_calculated
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_word_address_calculated
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_word_addrgen/$exit
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_word_addrgen/root_register_req
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_word_addrgen/root_register_ack
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_root_address_calculated
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_address_resized
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_word_addrgen/$entry
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_plus_offset/sum_rename_ack
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_complete/$exit
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_plus_offset/sum_rename_req
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_plus_offset/$exit
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/addr_of_3427_update_completed_
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_plus_offset/$entry
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_addr_resize/base_resize_ack
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_addr_resize/base_resize_req
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_addr_resize/$exit
      -- CP-element group 496: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_base_addr_resize/$entry
      -- 
    ack_7978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3427_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(496)); -- 
    -- CP-element group 497:  join  transition  output  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	490 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (9) 
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/ptr_deref_3430_Split/$exit
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/ptr_deref_3430_Split/$entry
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_sample_start_
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/ptr_deref_3430_Split/split_req
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/ptr_deref_3430_Split/split_ack
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/$entry
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/word_access_start/$entry
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/word_access_start/word_0/$entry
      -- CP-element group 497: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/word_access_start/word_0/rr
      -- 
    rr_8016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(497), ack => ptr_deref_3430_store_0_req_0); -- 
    zeropad3D_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(490) & zeropad3D_CP_2152_elements(496);
      gj_zeropad3D_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  transition  input  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498:  members (5) 
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_sample_completed_
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/$exit
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/word_access_start/$exit
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/word_access_start/word_0/$exit
      -- CP-element group 498: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Sample/word_access_start/word_0/ra
      -- 
    ra_8017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3430_store_0_ack_0, ack => zeropad3D_CP_2152_elements(498)); -- 
    -- CP-element group 499:  transition  input  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	465 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	500 
    -- CP-element group 499:  members (5) 
      -- CP-element group 499: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_update_completed_
      -- CP-element group 499: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/$exit
      -- CP-element group 499: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/word_access_complete/$exit
      -- CP-element group 499: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/word_access_complete/word_0/$exit
      -- CP-element group 499: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/ptr_deref_3430_Update/word_access_complete/word_0/ca
      -- 
    ca_8028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3430_store_0_ack_1, ack => zeropad3D_CP_2152_elements(499)); -- 
    -- CP-element group 500:  join  transition  place  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	485 
    -- CP-element group 500: 	493 
    -- CP-element group 500: 	499 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	1026 
    -- CP-element group 500:  members (5) 
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse956_ifx_xend1004
      -- CP-element group 500: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432__exit__
      -- CP-element group 500: 	 branch_block_stmt_714/assign_stmt_3332_to_assign_stmt_3432/$exit
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse956_ifx_xend1004_PhiReq/$entry
      -- CP-element group 500: 	 branch_block_stmt_714/ifx_xelse956_ifx_xend1004_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_500: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_500"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(485) & zeropad3D_CP_2152_elements(493) & zeropad3D_CP_2152_elements(499);
      gj_zeropad3D_cp_element_group_500 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(500), clk => clk, reset => reset); --
    end block;
    -- CP-element group 501:  transition  input  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	1026 
    -- CP-element group 501: successors 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Sample/ra
      -- 
    ra_8040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3438_inst_ack_0, ack => zeropad3D_CP_2152_elements(501)); -- 
    -- CP-element group 502:  branch  transition  place  input  output  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	1026 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502: 	504 
    -- CP-element group 502:  members (13) 
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452__exit__
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453__entry__
      -- CP-element group 502: 	 branch_block_stmt_714/R_cmp1012_3454_place
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/$exit
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_update_completed_
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Update/ca
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453_dead_link/$entry
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453_eval_test/$entry
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453_eval_test/$exit
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453_eval_test/branch_req
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453_if_link/$entry
      -- CP-element group 502: 	 branch_block_stmt_714/if_stmt_3453_else_link/$entry
      -- 
    ca_8045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3438_inst_ack_1, ack => zeropad3D_CP_2152_elements(502)); -- 
    branch_req_8053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(502), ack => if_stmt_3453_branch_req_0); -- 
    -- CP-element group 503:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	502 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	1035 
    -- CP-element group 503: 	1036 
    -- CP-element group 503: 	1038 
    -- CP-element group 503: 	1039 
    -- CP-element group 503: 	1041 
    -- CP-element group 503: 	1042 
    -- CP-element group 503:  members (40) 
      -- CP-element group 503: 	 branch_block_stmt_714/merge_stmt_3459__exit__
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3465__exit__
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3465__entry__
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xend1004_ifx_xthen1014
      -- CP-element group 503: 	 branch_block_stmt_714/if_stmt_3453_if_link/$exit
      -- CP-element group 503: 	 branch_block_stmt_714/if_stmt_3453_if_link/if_choice_transition
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3465/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/assign_stmt_3465/$exit
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xend1004_ifx_xthen1014_PhiReq/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xend1004_ifx_xthen1014_PhiReq/$exit
      -- CP-element group 503: 	 branch_block_stmt_714/merge_stmt_3459_PhiReqMerge
      -- CP-element group 503: 	 branch_block_stmt_714/merge_stmt_3459_PhiAck/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/merge_stmt_3459_PhiAck/$exit
      -- CP-element group 503: 	 branch_block_stmt_714/merge_stmt_3459_PhiAck/dummy
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Sample/rr
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Update/cr
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Sample/rr
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Update/cr
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Sample/rr
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3453_branch_ack_1, ack => zeropad3D_CP_2152_elements(503)); -- 
    rr_13255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(503), ack => type_cast_3562_inst_req_0); -- 
    cr_13260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(503), ack => type_cast_3562_inst_req_1); -- 
    rr_13278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(503), ack => type_cast_3569_inst_req_0); -- 
    cr_13283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(503), ack => type_cast_3569_inst_req_1); -- 
    rr_13301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(503), ack => type_cast_3577_inst_req_0); -- 
    cr_13306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(503), ack => type_cast_3577_inst_req_1); -- 
    -- CP-element group 504:  fork  transition  place  input  output  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	502 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	505 
    -- CP-element group 504: 	506 
    -- CP-element group 504: 	507 
    -- CP-element group 504: 	508 
    -- CP-element group 504: 	510 
    -- CP-element group 504: 	513 
    -- CP-element group 504: 	515 
    -- CP-element group 504: 	516 
    -- CP-element group 504: 	517 
    -- CP-element group 504: 	519 
    -- CP-element group 504:  members (54) 
      -- CP-element group 504: 	 branch_block_stmt_714/merge_stmt_3467__exit__
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551__entry__
      -- CP-element group 504: 	 branch_block_stmt_714/ifx_xend1004_ifx_xelse1019
      -- CP-element group 504: 	 branch_block_stmt_714/if_stmt_3453_else_link/$exit
      -- CP-element group 504: 	 branch_block_stmt_714/if_stmt_3453_else_link/else_choice_transition
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_sample_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Sample/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Sample/rr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_sample_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_word_address_calculated
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_root_address_calculated
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/word_access_start/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/word_access_start/word_0/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/word_access_start/word_0/rr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/word_access_complete/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/word_access_complete/word_0/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/word_access_complete/word_0/cr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_sample_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_word_address_calculated
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_root_address_calculated
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/word_access_start/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/word_access_start/word_0/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/word_access_start/word_0/rr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/word_access_complete/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/word_access_complete/word_0/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/word_access_complete/word_0/cr
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_update_start_
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_714/ifx_xend1004_ifx_xelse1019_PhiReq/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/ifx_xend1004_ifx_xelse1019_PhiReq/$exit
      -- CP-element group 504: 	 branch_block_stmt_714/merge_stmt_3467_PhiReqMerge
      -- CP-element group 504: 	 branch_block_stmt_714/merge_stmt_3467_PhiAck/$entry
      -- CP-element group 504: 	 branch_block_stmt_714/merge_stmt_3467_PhiAck/$exit
      -- CP-element group 504: 	 branch_block_stmt_714/merge_stmt_3467_PhiAck/dummy
      -- 
    else_choice_transition_8062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3453_branch_ack_0, ack => zeropad3D_CP_2152_elements(504)); -- 
    rr_8078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => type_cast_3477_inst_req_0); -- 
    cr_8083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => type_cast_3477_inst_req_1); -- 
    rr_8100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => LOAD_col_high_3480_load_0_req_0); -- 
    cr_8111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => LOAD_col_high_3480_load_0_req_1); -- 
    cr_8130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => type_cast_3484_inst_req_1); -- 
    cr_8144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => type_cast_3504_inst_req_1); -- 
    cr_8158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => type_cast_3521_inst_req_1); -- 
    rr_8175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => LOAD_row_high_3524_load_0_req_0); -- 
    cr_8186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => LOAD_row_high_3524_load_0_req_1); -- 
    cr_8205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(504), ack => type_cast_3528_inst_req_1); -- 
    -- CP-element group 505:  transition  input  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	504 
    -- CP-element group 505: successors 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_sample_completed_
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Sample/$exit
      -- CP-element group 505: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Sample/ra
      -- 
    ra_8079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3477_inst_ack_0, ack => zeropad3D_CP_2152_elements(505)); -- 
    -- CP-element group 506:  transition  input  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	504 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	511 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_update_completed_
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Update/$exit
      -- CP-element group 506: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3477_Update/ca
      -- 
    ca_8084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3477_inst_ack_1, ack => zeropad3D_CP_2152_elements(506)); -- 
    -- CP-element group 507:  transition  input  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	504 
    -- CP-element group 507: successors 
    -- CP-element group 507:  members (5) 
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_sample_completed_
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/$exit
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/word_access_start/$exit
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/word_access_start/word_0/$exit
      -- CP-element group 507: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Sample/word_access_start/word_0/ra
      -- 
    ra_8101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3480_load_0_ack_0, ack => zeropad3D_CP_2152_elements(507)); -- 
    -- CP-element group 508:  transition  input  output  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	504 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	509 
    -- CP-element group 508:  members (12) 
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_update_completed_
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/word_access_complete/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/word_access_complete/word_0/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/word_access_complete/word_0/ca
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/LOAD_col_high_3480_Merge/$entry
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/LOAD_col_high_3480_Merge/$exit
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/LOAD_col_high_3480_Merge/merge_req
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_col_high_3480_Update/LOAD_col_high_3480_Merge/merge_ack
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_sample_start_
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Sample/$entry
      -- CP-element group 508: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Sample/rr
      -- 
    ca_8112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3480_load_0_ack_1, ack => zeropad3D_CP_2152_elements(508)); -- 
    rr_8125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(508), ack => type_cast_3484_inst_req_0); -- 
    -- CP-element group 509:  transition  input  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	508 
    -- CP-element group 509: successors 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_sample_completed_
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Sample/$exit
      -- CP-element group 509: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Sample/ra
      -- 
    ra_8126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3484_inst_ack_0, ack => zeropad3D_CP_2152_elements(509)); -- 
    -- CP-element group 510:  transition  input  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	504 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	511 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_update_completed_
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Update/$exit
      -- CP-element group 510: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3484_Update/ca
      -- 
    ca_8131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3484_inst_ack_1, ack => zeropad3D_CP_2152_elements(510)); -- 
    -- CP-element group 511:  join  transition  output  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	506 
    -- CP-element group 511: 	510 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	512 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_sample_start_
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Sample/$entry
      -- CP-element group 511: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Sample/rr
      -- 
    rr_8139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(511), ack => type_cast_3504_inst_req_0); -- 
    zeropad3D_cp_element_group_511: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_511"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(506) & zeropad3D_CP_2152_elements(510);
      gj_zeropad3D_cp_element_group_511 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(511), clk => clk, reset => reset); --
    end block;
    -- CP-element group 512:  transition  input  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	511 
    -- CP-element group 512: successors 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_sample_completed_
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Sample/$exit
      -- CP-element group 512: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Sample/ra
      -- 
    ra_8140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3504_inst_ack_0, ack => zeropad3D_CP_2152_elements(512)); -- 
    -- CP-element group 513:  transition  input  output  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	504 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	514 
    -- CP-element group 513:  members (6) 
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_update_completed_
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Update/$exit
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3504_Update/ca
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_sample_start_
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Sample/$entry
      -- CP-element group 513: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Sample/rr
      -- 
    ca_8145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3504_inst_ack_1, ack => zeropad3D_CP_2152_elements(513)); -- 
    rr_8153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(513), ack => type_cast_3521_inst_req_0); -- 
    -- CP-element group 514:  transition  input  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	513 
    -- CP-element group 514: successors 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_sample_completed_
      -- CP-element group 514: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Sample/$exit
      -- CP-element group 514: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Sample/ra
      -- 
    ra_8154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3521_inst_ack_0, ack => zeropad3D_CP_2152_elements(514)); -- 
    -- CP-element group 515:  transition  input  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	504 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	520 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_update_completed_
      -- CP-element group 515: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Update/$exit
      -- CP-element group 515: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3521_Update/ca
      -- 
    ca_8159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 515_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3521_inst_ack_1, ack => zeropad3D_CP_2152_elements(515)); -- 
    -- CP-element group 516:  transition  input  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	504 
    -- CP-element group 516: successors 
    -- CP-element group 516:  members (5) 
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_sample_completed_
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/$exit
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/word_access_start/$exit
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/word_access_start/word_0/$exit
      -- CP-element group 516: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Sample/word_access_start/word_0/ra
      -- 
    ra_8176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3524_load_0_ack_0, ack => zeropad3D_CP_2152_elements(516)); -- 
    -- CP-element group 517:  transition  input  output  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	504 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	518 
    -- CP-element group 517:  members (12) 
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_update_completed_
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/$exit
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/word_access_complete/$exit
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/word_access_complete/word_0/$exit
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/word_access_complete/word_0/ca
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/LOAD_row_high_3524_Merge/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/LOAD_row_high_3524_Merge/$exit
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/LOAD_row_high_3524_Merge/merge_req
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/LOAD_row_high_3524_Update/LOAD_row_high_3524_Merge/merge_ack
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_sample_start_
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Sample/$entry
      -- CP-element group 517: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Sample/rr
      -- 
    ca_8187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3524_load_0_ack_1, ack => zeropad3D_CP_2152_elements(517)); -- 
    rr_8200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(517), ack => type_cast_3528_inst_req_0); -- 
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	517 
    -- CP-element group 518: successors 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_sample_completed_
      -- CP-element group 518: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Sample/$exit
      -- CP-element group 518: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Sample/ra
      -- 
    ra_8201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3528_inst_ack_0, ack => zeropad3D_CP_2152_elements(518)); -- 
    -- CP-element group 519:  transition  input  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	504 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	520 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_update_completed_
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Update/$exit
      -- CP-element group 519: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/type_cast_3528_Update/ca
      -- 
    ca_8206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3528_inst_ack_1, ack => zeropad3D_CP_2152_elements(519)); -- 
    -- CP-element group 520:  branch  join  transition  place  output  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	515 
    -- CP-element group 520: 	519 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	521 
    -- CP-element group 520: 	522 
    -- CP-element group 520:  members (10) 
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552__entry__
      -- CP-element group 520: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551__exit__
      -- CP-element group 520: 	 branch_block_stmt_714/R_cmp1048_3553_place
      -- CP-element group 520: 	 branch_block_stmt_714/assign_stmt_3473_to_assign_stmt_3551/$exit
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552_dead_link/$entry
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552_eval_test/$entry
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552_eval_test/$exit
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552_eval_test/branch_req
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552_if_link/$entry
      -- CP-element group 520: 	 branch_block_stmt_714/if_stmt_3552_else_link/$entry
      -- 
    branch_req_8214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(520), ack => if_stmt_3552_branch_req_0); -- 
    zeropad3D_cp_element_group_520: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_520"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(515) & zeropad3D_CP_2152_elements(519);
      gj_zeropad3D_cp_element_group_520 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(520), clk => clk, reset => reset); --
    end block;
    -- CP-element group 521:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	520 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	523 
    -- CP-element group 521: 	524 
    -- CP-element group 521: 	526 
    -- CP-element group 521: 	527 
    -- CP-element group 521: 	528 
    -- CP-element group 521: 	530 
    -- CP-element group 521: 	531 
    -- CP-element group 521: 	532 
    -- CP-element group 521: 	533 
    -- CP-element group 521: 	534 
    -- CP-element group 521: 	535 
    -- CP-element group 521: 	536 
    -- CP-element group 521: 	537 
    -- CP-element group 521: 	538 
    -- CP-element group 521: 	540 
    -- CP-element group 521: 	542 
    -- CP-element group 521: 	544 
    -- CP-element group 521:  members (127) 
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725__entry__
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3580__exit__
      -- CP-element group 521: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058
      -- CP-element group 521: 	 branch_block_stmt_714/if_stmt_3552_if_link/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/if_stmt_3552_if_link/if_choice_transition
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_address_resized
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_addr_resize/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_addr_resize/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_addr_resize/base_resize_req
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_addr_resize/base_resize_ack
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_plus_offset/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_plus_offset/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_plus_offset/sum_rename_req
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_base_plus_offset/sum_rename_ack
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_word_addrgen/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_word_addrgen/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_word_addrgen/root_register_req
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_word_addrgen/root_register_ack
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_sample_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_word_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_root_address_calculated
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_address_resized
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_addr_resize/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_addr_resize/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_addr_resize/base_resize_req
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_addr_resize/base_resize_ack
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_plus_offset/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_plus_offset/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_plus_offset/sum_rename_req
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_base_plus_offset/sum_rename_ack
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_word_addrgen/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_word_addrgen/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_word_addrgen/root_register_req
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_word_addrgen/root_register_ack
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/word_access_start/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/word_access_start/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/word_access_start/word_0/rr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_update_start_
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/ifx_xelse1019_whilex_xend1058_PhiReq/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3580_PhiReqMerge
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3580_PhiAck/$entry
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3580_PhiAck/$exit
      -- CP-element group 521: 	 branch_block_stmt_714/merge_stmt_3580_PhiAck/dummy
      -- 
    if_choice_transition_8219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3552_branch_ack_1, ack => zeropad3D_CP_2152_elements(521)); -- 
    rr_8244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_col_high_3583_load_0_req_0); -- 
    cr_8255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_col_high_3583_load_0_req_1); -- 
    cr_8274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => type_cast_3587_inst_req_1); -- 
    rr_8291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_row_high_3596_load_0_req_0); -- 
    cr_8302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_row_high_3596_load_0_req_1); -- 
    cr_8321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => type_cast_3600_inst_req_1); -- 
    rr_8338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_pad_3609_load_0_req_0); -- 
    cr_8349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_pad_3609_load_0_req_1); -- 
    rr_8371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_depth_high_3612_load_0_req_0); -- 
    cr_8382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => LOAD_depth_high_3612_load_0_req_1); -- 
    rr_8421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => ptr_deref_3624_load_0_req_0); -- 
    cr_8432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => ptr_deref_3624_load_0_req_1); -- 
    rr_8471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => ptr_deref_3636_load_0_req_0); -- 
    cr_8482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => ptr_deref_3636_load_0_req_1); -- 
    cr_8501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => type_cast_3640_inst_req_1); -- 
    cr_8515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => type_cast_3644_inst_req_1); -- 
    cr_8529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(521), ack => type_cast_3683_inst_req_1); -- 
    -- CP-element group 522:  fork  transition  place  input  output  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	520 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	1027 
    -- CP-element group 522: 	1028 
    -- CP-element group 522: 	1029 
    -- CP-element group 522: 	1031 
    -- CP-element group 522: 	1032 
    -- CP-element group 522:  members (22) 
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057
      -- CP-element group 522: 	 branch_block_stmt_714/if_stmt_3552_else_link/$exit
      -- CP-element group 522: 	 branch_block_stmt_714/if_stmt_3552_else_link/else_choice_transition
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3559/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Sample/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Sample/rr
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Update/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Update/cr
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Sample/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Sample/rr
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Update/$entry
      -- CP-element group 522: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3552_branch_ack_0, ack => zeropad3D_CP_2152_elements(522)); -- 
    rr_13206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(522), ack => type_cast_3571_inst_req_0); -- 
    cr_13211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(522), ack => type_cast_3571_inst_req_1); -- 
    rr_13229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(522), ack => type_cast_3575_inst_req_0); -- 
    cr_13234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(522), ack => type_cast_3575_inst_req_1); -- 
    -- CP-element group 523:  transition  input  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	521 
    -- CP-element group 523: successors 
    -- CP-element group 523:  members (5) 
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_sample_completed_
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/word_access_start/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/word_access_start/word_0/$exit
      -- CP-element group 523: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Sample/word_access_start/word_0/ra
      -- 
    ra_8245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3583_load_0_ack_0, ack => zeropad3D_CP_2152_elements(523)); -- 
    -- CP-element group 524:  fork  transition  input  output  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	521 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	525 
    -- CP-element group 524: 	541 
    -- CP-element group 524:  members (15) 
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_update_completed_
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/$exit
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/word_access_complete/$exit
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/word_access_complete/word_0/$exit
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/word_access_complete/word_0/ca
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/LOAD_col_high_3583_Merge/$entry
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/LOAD_col_high_3583_Merge/$exit
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/LOAD_col_high_3583_Merge/merge_req
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_col_high_3583_Update/LOAD_col_high_3583_Merge/merge_ack
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_sample_start_
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Sample/$entry
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Sample/rr
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_sample_start_
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Sample/$entry
      -- CP-element group 524: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Sample/rr
      -- 
    ca_8256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3583_load_0_ack_1, ack => zeropad3D_CP_2152_elements(524)); -- 
    rr_8269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(524), ack => type_cast_3587_inst_req_0); -- 
    rr_8510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(524), ack => type_cast_3644_inst_req_0); -- 
    -- CP-element group 525:  transition  input  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	524 
    -- CP-element group 525: successors 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_sample_completed_
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Sample/$exit
      -- CP-element group 525: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Sample/ra
      -- 
    ra_8270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3587_inst_ack_0, ack => zeropad3D_CP_2152_elements(525)); -- 
    -- CP-element group 526:  transition  input  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	521 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	545 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_update_completed_
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Update/$exit
      -- CP-element group 526: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3587_Update/ca
      -- 
    ca_8275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 526_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3587_inst_ack_1, ack => zeropad3D_CP_2152_elements(526)); -- 
    -- CP-element group 527:  transition  input  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	521 
    -- CP-element group 527: successors 
    -- CP-element group 527:  members (5) 
      -- CP-element group 527: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_sample_completed_
      -- CP-element group 527: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/$exit
      -- CP-element group 527: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/word_access_start/$exit
      -- CP-element group 527: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/word_access_start/word_0/$exit
      -- CP-element group 527: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Sample/word_access_start/word_0/ra
      -- 
    ra_8292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3596_load_0_ack_0, ack => zeropad3D_CP_2152_elements(527)); -- 
    -- CP-element group 528:  transition  input  output  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	521 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	529 
    -- CP-element group 528:  members (12) 
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_update_completed_
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/$exit
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/word_access_complete/$exit
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/word_access_complete/word_0/$exit
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/word_access_complete/word_0/ca
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/LOAD_row_high_3596_Merge/$entry
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/LOAD_row_high_3596_Merge/$exit
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/LOAD_row_high_3596_Merge/merge_req
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_row_high_3596_Update/LOAD_row_high_3596_Merge/merge_ack
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Sample/rr
      -- 
    ca_8303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3596_load_0_ack_1, ack => zeropad3D_CP_2152_elements(528)); -- 
    rr_8316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(528), ack => type_cast_3600_inst_req_0); -- 
    -- CP-element group 529:  transition  input  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	528 
    -- CP-element group 529: successors 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_sample_completed_
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Sample/$exit
      -- CP-element group 529: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Sample/ra
      -- 
    ra_8317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 529_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3600_inst_ack_0, ack => zeropad3D_CP_2152_elements(529)); -- 
    -- CP-element group 530:  transition  input  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	521 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	545 
    -- CP-element group 530:  members (3) 
      -- CP-element group 530: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_update_completed_
      -- CP-element group 530: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Update/$exit
      -- CP-element group 530: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3600_Update/ca
      -- 
    ca_8322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3600_inst_ack_1, ack => zeropad3D_CP_2152_elements(530)); -- 
    -- CP-element group 531:  transition  input  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	521 
    -- CP-element group 531: successors 
    -- CP-element group 531:  members (5) 
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_sample_completed_
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/$exit
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/word_access_start/$exit
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/word_access_start/word_0/$exit
      -- CP-element group 531: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Sample/word_access_start/word_0/ra
      -- 
    ra_8339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3609_load_0_ack_0, ack => zeropad3D_CP_2152_elements(531)); -- 
    -- CP-element group 532:  transition  input  output  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	521 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	543 
    -- CP-element group 532:  members (12) 
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_update_completed_
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/word_access_complete/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/word_access_complete/word_0/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/word_access_complete/word_0/ca
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/LOAD_pad_3609_Merge/$entry
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/LOAD_pad_3609_Merge/$exit
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/LOAD_pad_3609_Merge/merge_req
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_pad_3609_Update/LOAD_pad_3609_Merge/merge_ack
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_sample_start_
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Sample/$entry
      -- CP-element group 532: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Sample/rr
      -- 
    ca_8350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3609_load_0_ack_1, ack => zeropad3D_CP_2152_elements(532)); -- 
    rr_8524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(532), ack => type_cast_3683_inst_req_0); -- 
    -- CP-element group 533:  transition  input  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	521 
    -- CP-element group 533: successors 
    -- CP-element group 533:  members (5) 
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_sample_completed_
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/word_access_start/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/word_access_start/word_0/$exit
      -- CP-element group 533: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Sample/word_access_start/word_0/ra
      -- 
    ra_8372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3612_load_0_ack_0, ack => zeropad3D_CP_2152_elements(533)); -- 
    -- CP-element group 534:  transition  input  output  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	521 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	539 
    -- CP-element group 534:  members (12) 
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_update_completed_
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/$exit
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/word_access_complete/$exit
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/word_access_complete/word_0/$exit
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/word_access_complete/word_0/ca
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/LOAD_depth_high_3612_Merge/$entry
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/LOAD_depth_high_3612_Merge/$exit
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/LOAD_depth_high_3612_Merge/merge_req
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/LOAD_depth_high_3612_Update/LOAD_depth_high_3612_Merge/merge_ack
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_sample_start_
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Sample/$entry
      -- CP-element group 534: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Sample/rr
      -- 
    ca_8383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_3612_load_0_ack_1, ack => zeropad3D_CP_2152_elements(534)); -- 
    rr_8496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(534), ack => type_cast_3640_inst_req_0); -- 
    -- CP-element group 535:  transition  input  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	521 
    -- CP-element group 535: successors 
    -- CP-element group 535:  members (5) 
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_sample_completed_
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/$exit
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/word_access_start/$exit
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/word_access_start/word_0/$exit
      -- CP-element group 535: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Sample/word_access_start/word_0/ra
      -- 
    ra_8422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3624_load_0_ack_0, ack => zeropad3D_CP_2152_elements(535)); -- 
    -- CP-element group 536:  transition  input  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	521 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	545 
    -- CP-element group 536:  members (9) 
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_update_completed_
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/word_access_complete/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/word_access_complete/word_0/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/word_access_complete/word_0/ca
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/ptr_deref_3624_Merge/$entry
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/ptr_deref_3624_Merge/$exit
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/ptr_deref_3624_Merge/merge_req
      -- CP-element group 536: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3624_Update/ptr_deref_3624_Merge/merge_ack
      -- 
    ca_8433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3624_load_0_ack_1, ack => zeropad3D_CP_2152_elements(536)); -- 
    -- CP-element group 537:  transition  input  bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	521 
    -- CP-element group 537: successors 
    -- CP-element group 537:  members (5) 
      -- CP-element group 537: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_sample_completed_
      -- CP-element group 537: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/$exit
      -- CP-element group 537: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/word_access_start/$exit
      -- CP-element group 537: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/word_access_start/word_0/$exit
      -- CP-element group 537: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Sample/word_access_start/word_0/ra
      -- 
    ra_8472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3636_load_0_ack_0, ack => zeropad3D_CP_2152_elements(537)); -- 
    -- CP-element group 538:  transition  input  bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	521 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	545 
    -- CP-element group 538:  members (9) 
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_update_completed_
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/$exit
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/word_access_complete/$exit
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/word_access_complete/word_0/$exit
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/word_access_complete/word_0/ca
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/ptr_deref_3636_Merge/$entry
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/ptr_deref_3636_Merge/$exit
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/ptr_deref_3636_Merge/merge_req
      -- CP-element group 538: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/ptr_deref_3636_Update/ptr_deref_3636_Merge/merge_ack
      -- 
    ca_8483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 538_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3636_load_0_ack_1, ack => zeropad3D_CP_2152_elements(538)); -- 
    -- CP-element group 539:  transition  input  bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	534 
    -- CP-element group 539: successors 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_sample_completed_
      -- CP-element group 539: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Sample/ra
      -- 
    ra_8497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3640_inst_ack_0, ack => zeropad3D_CP_2152_elements(539)); -- 
    -- CP-element group 540:  transition  input  bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	521 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	545 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_update_completed_
      -- CP-element group 540: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3640_Update/ca
      -- 
    ca_8502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3640_inst_ack_1, ack => zeropad3D_CP_2152_elements(540)); -- 
    -- CP-element group 541:  transition  input  bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	524 
    -- CP-element group 541: successors 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_sample_completed_
      -- CP-element group 541: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Sample/$exit
      -- CP-element group 541: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Sample/ra
      -- 
    ra_8511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3644_inst_ack_0, ack => zeropad3D_CP_2152_elements(541)); -- 
    -- CP-element group 542:  transition  input  bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	521 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	545 
    -- CP-element group 542:  members (3) 
      -- CP-element group 542: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_update_completed_
      -- CP-element group 542: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Update/$exit
      -- CP-element group 542: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3644_Update/ca
      -- 
    ca_8516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3644_inst_ack_1, ack => zeropad3D_CP_2152_elements(542)); -- 
    -- CP-element group 543:  transition  input  bypass 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	532 
    -- CP-element group 543: successors 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_sample_completed_
      -- CP-element group 543: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Sample/$exit
      -- CP-element group 543: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Sample/ra
      -- 
    ra_8525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3683_inst_ack_0, ack => zeropad3D_CP_2152_elements(543)); -- 
    -- CP-element group 544:  transition  input  bypass 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	521 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	545 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_update_completed_
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Update/$exit
      -- CP-element group 544: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/type_cast_3683_Update/ca
      -- 
    ca_8530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3683_inst_ack_1, ack => zeropad3D_CP_2152_elements(544)); -- 
    -- CP-element group 545:  join  fork  transition  place  output  bypass 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	526 
    -- CP-element group 545: 	530 
    -- CP-element group 545: 	536 
    -- CP-element group 545: 	538 
    -- CP-element group 545: 	540 
    -- CP-element group 545: 	542 
    -- CP-element group 545: 	544 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	1060 
    -- CP-element group 545: 	1061 
    -- CP-element group 545: 	1062 
    -- CP-element group 545: 	1064 
    -- CP-element group 545: 	1065 
    -- CP-element group 545:  members (22) 
      -- CP-element group 545: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725__exit__
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122
      -- CP-element group 545: 	 branch_block_stmt_714/assign_stmt_3584_to_assign_stmt_3725/$exit
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3728/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Sample/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Sample/rr
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Update/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Update/cr
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Sample/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Sample/rr
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Update/$entry
      -- CP-element group 545: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Update/cr
      -- 
    rr_13422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(545), ack => type_cast_3738_inst_req_0); -- 
    cr_13427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(545), ack => type_cast_3738_inst_req_1); -- 
    rr_13445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(545), ack => type_cast_3746_inst_req_0); -- 
    cr_13450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(545), ack => type_cast_3746_inst_req_1); -- 
    zeropad3D_cp_element_group_545: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_545"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(526) & zeropad3D_CP_2152_elements(530) & zeropad3D_CP_2152_elements(536) & zeropad3D_CP_2152_elements(538) & zeropad3D_CP_2152_elements(540) & zeropad3D_CP_2152_elements(542) & zeropad3D_CP_2152_elements(544);
      gj_zeropad3D_cp_element_group_545 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(545), clk => clk, reset => reset); --
    end block;
    -- CP-element group 546:  transition  input  bypass 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	1072 
    -- CP-element group 546: successors 
    -- CP-element group 546:  members (3) 
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_sample_completed_
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Sample/$exit
      -- CP-element group 546: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Sample/ra
      -- 
    ra_8542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3751_inst_ack_0, ack => zeropad3D_CP_2152_elements(546)); -- 
    -- CP-element group 547:  branch  transition  place  input  output  bypass 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	1072 
    -- CP-element group 547: successors 
    -- CP-element group 547: 	548 
    -- CP-element group 547: 	549 
    -- CP-element group 547:  members (13) 
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759__exit__
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760__entry__
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/$exit
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_update_completed_
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Update/$exit
      -- CP-element group 547: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Update/ca
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760_dead_link/$entry
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760_eval_test/$entry
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760_eval_test/$exit
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760_eval_test/branch_req
      -- CP-element group 547: 	 branch_block_stmt_714/R_cmp1127_3761_place
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760_if_link/$entry
      -- CP-element group 547: 	 branch_block_stmt_714/if_stmt_3760_else_link/$entry
      -- 
    ca_8547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3751_inst_ack_1, ack => zeropad3D_CP_2152_elements(547)); -- 
    branch_req_8555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(547), ack => if_stmt_3760_branch_req_0); -- 
    -- CP-element group 548:  transition  place  input  bypass 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	547 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	1073 
    -- CP-element group 548:  members (5) 
      -- CP-element group 548: 	 branch_block_stmt_714/if_stmt_3760_if_link/$exit
      -- CP-element group 548: 	 branch_block_stmt_714/if_stmt_3760_if_link/if_choice_transition
      -- CP-element group 548: 	 branch_block_stmt_714/whilex_xbody1122_ifx_xthen1158
      -- CP-element group 548: 	 branch_block_stmt_714/whilex_xbody1122_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 548: 	 branch_block_stmt_714/whilex_xbody1122_ifx_xthen1158_PhiReq/$exit
      -- 
    if_choice_transition_8560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3760_branch_ack_1, ack => zeropad3D_CP_2152_elements(548)); -- 
    -- CP-element group 549:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	547 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	550 
    -- CP-element group 549: 	551 
    -- CP-element group 549: 	553 
    -- CP-element group 549:  members (27) 
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797__entry__
      -- CP-element group 549: 	 branch_block_stmt_714/merge_stmt_3766__exit__
      -- CP-element group 549: 	 branch_block_stmt_714/if_stmt_3760_else_link/$exit
      -- CP-element group 549: 	 branch_block_stmt_714/if_stmt_3760_else_link/else_choice_transition
      -- CP-element group 549: 	 branch_block_stmt_714/whilex_xbody1122_lorx_xlhsx_xfalse1129
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_sample_start_
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_update_start_
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_word_address_calculated
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_root_address_calculated
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/word_access_start/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/word_access_start/word_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/word_access_start/word_0/rr
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/word_access_complete/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/word_access_complete/word_0/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/word_access_complete/word_0/cr
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_update_start_
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Update/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Update/cr
      -- CP-element group 549: 	 branch_block_stmt_714/whilex_xbody1122_lorx_xlhsx_xfalse1129_PhiReq/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/whilex_xbody1122_lorx_xlhsx_xfalse1129_PhiReq/$exit
      -- CP-element group 549: 	 branch_block_stmt_714/merge_stmt_3766_PhiReqMerge
      -- CP-element group 549: 	 branch_block_stmt_714/merge_stmt_3766_PhiAck/$entry
      -- CP-element group 549: 	 branch_block_stmt_714/merge_stmt_3766_PhiAck/$exit
      -- CP-element group 549: 	 branch_block_stmt_714/merge_stmt_3766_PhiAck/dummy
      -- 
    else_choice_transition_8564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3760_branch_ack_0, ack => zeropad3D_CP_2152_elements(549)); -- 
    rr_8585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(549), ack => LOAD_row_high_3768_load_0_req_0); -- 
    cr_8596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(549), ack => LOAD_row_high_3768_load_0_req_1); -- 
    cr_8615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(549), ack => type_cast_3772_inst_req_1); -- 
    -- CP-element group 550:  transition  input  bypass 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	549 
    -- CP-element group 550: successors 
    -- CP-element group 550:  members (5) 
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_sample_completed_
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/$exit
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/word_access_start/$exit
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/word_access_start/word_0/$exit
      -- CP-element group 550: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Sample/word_access_start/word_0/ra
      -- 
    ra_8586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3768_load_0_ack_0, ack => zeropad3D_CP_2152_elements(550)); -- 
    -- CP-element group 551:  transition  input  output  bypass 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	549 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	552 
    -- CP-element group 551:  members (12) 
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_update_completed_
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/$exit
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/word_access_complete/$exit
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/word_access_complete/word_0/$exit
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/word_access_complete/word_0/ca
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/LOAD_row_high_3768_Merge/$entry
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/LOAD_row_high_3768_Merge/$exit
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/LOAD_row_high_3768_Merge/merge_req
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/LOAD_row_high_3768_Update/LOAD_row_high_3768_Merge/merge_ack
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_sample_start_
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Sample/$entry
      -- CP-element group 551: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Sample/rr
      -- 
    ca_8597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 551_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_3768_load_0_ack_1, ack => zeropad3D_CP_2152_elements(551)); -- 
    rr_8610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(551), ack => type_cast_3772_inst_req_0); -- 
    -- CP-element group 552:  transition  input  bypass 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	551 
    -- CP-element group 552: successors 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_sample_completed_
      -- CP-element group 552: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Sample/$exit
      -- CP-element group 552: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Sample/ra
      -- 
    ra_8611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3772_inst_ack_0, ack => zeropad3D_CP_2152_elements(552)); -- 
    -- CP-element group 553:  branch  transition  place  input  output  bypass 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	549 
    -- CP-element group 553: successors 
    -- CP-element group 553: 	554 
    -- CP-element group 553: 	555 
    -- CP-element group 553:  members (13) 
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797__exit__
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798__entry__
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/$exit
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Update/$exit
      -- CP-element group 553: 	 branch_block_stmt_714/assign_stmt_3769_to_assign_stmt_3797/type_cast_3772_Update/ca
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798_dead_link/$entry
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798_eval_test/$entry
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798_eval_test/$exit
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798_eval_test/branch_req
      -- CP-element group 553: 	 branch_block_stmt_714/R_cmp1139_3799_place
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798_if_link/$entry
      -- CP-element group 553: 	 branch_block_stmt_714/if_stmt_3798_else_link/$entry
      -- 
    ca_8616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3772_inst_ack_1, ack => zeropad3D_CP_2152_elements(553)); -- 
    branch_req_8624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(553), ack => if_stmt_3798_branch_req_0); -- 
    -- CP-element group 554:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	553 
    -- CP-element group 554: successors 
    -- CP-element group 554: 	556 
    -- CP-element group 554: 	557 
    -- CP-element group 554:  members (18) 
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816__entry__
      -- CP-element group 554: 	 branch_block_stmt_714/merge_stmt_3804__exit__
      -- CP-element group 554: 	 branch_block_stmt_714/if_stmt_3798_if_link/$exit
      -- CP-element group 554: 	 branch_block_stmt_714/if_stmt_3798_if_link/if_choice_transition
      -- CP-element group 554: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_lorx_xlhsx_xfalse1141
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/$entry
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_sample_start_
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_update_start_
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Sample/$entry
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Sample/rr
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Update/$entry
      -- CP-element group 554: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Update/cr
      -- CP-element group 554: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_lorx_xlhsx_xfalse1141_PhiReq/$entry
      -- CP-element group 554: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_lorx_xlhsx_xfalse1141_PhiReq/$exit
      -- CP-element group 554: 	 branch_block_stmt_714/merge_stmt_3804_PhiReqMerge
      -- CP-element group 554: 	 branch_block_stmt_714/merge_stmt_3804_PhiAck/$entry
      -- CP-element group 554: 	 branch_block_stmt_714/merge_stmt_3804_PhiAck/$exit
      -- CP-element group 554: 	 branch_block_stmt_714/merge_stmt_3804_PhiAck/dummy
      -- 
    if_choice_transition_8629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 554_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3798_branch_ack_1, ack => zeropad3D_CP_2152_elements(554)); -- 
    rr_8646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(554), ack => type_cast_3808_inst_req_0); -- 
    cr_8651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(554), ack => type_cast_3808_inst_req_1); -- 
    -- CP-element group 555:  transition  place  input  bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	553 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	1073 
    -- CP-element group 555:  members (5) 
      -- CP-element group 555: 	 branch_block_stmt_714/if_stmt_3798_else_link/$exit
      -- CP-element group 555: 	 branch_block_stmt_714/if_stmt_3798_else_link/else_choice_transition
      -- CP-element group 555: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_ifx_xthen1158
      -- CP-element group 555: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 555: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1129_ifx_xthen1158_PhiReq/$exit
      -- 
    else_choice_transition_8633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 555_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3798_branch_ack_0, ack => zeropad3D_CP_2152_elements(555)); -- 
    -- CP-element group 556:  transition  input  bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	554 
    -- CP-element group 556: successors 
    -- CP-element group 556:  members (3) 
      -- CP-element group 556: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_sample_completed_
      -- CP-element group 556: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Sample/$exit
      -- CP-element group 556: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Sample/ra
      -- 
    ra_8647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3808_inst_ack_0, ack => zeropad3D_CP_2152_elements(556)); -- 
    -- CP-element group 557:  branch  transition  place  input  output  bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	554 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	558 
    -- CP-element group 557: 	559 
    -- CP-element group 557:  members (13) 
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816__exit__
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817__entry__
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/$exit
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_update_completed_
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Update/$exit
      -- CP-element group 557: 	 branch_block_stmt_714/assign_stmt_3809_to_assign_stmt_3816/type_cast_3808_Update/ca
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817_dead_link/$entry
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817_eval_test/$entry
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817_eval_test/$exit
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817_eval_test/branch_req
      -- CP-element group 557: 	 branch_block_stmt_714/R_cmp1146_3818_place
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817_if_link/$entry
      -- CP-element group 557: 	 branch_block_stmt_714/if_stmt_3817_else_link/$entry
      -- 
    ca_8652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3808_inst_ack_1, ack => zeropad3D_CP_2152_elements(557)); -- 
    branch_req_8660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(557), ack => if_stmt_3817_branch_req_0); -- 
    -- CP-element group 558:  transition  place  input  bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	557 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	1073 
    -- CP-element group 558:  members (5) 
      -- CP-element group 558: 	 branch_block_stmt_714/if_stmt_3817_if_link/$exit
      -- CP-element group 558: 	 branch_block_stmt_714/if_stmt_3817_if_link/if_choice_transition
      -- CP-element group 558: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_ifx_xthen1158
      -- CP-element group 558: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 558: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_ifx_xthen1158_PhiReq/$exit
      -- 
    if_choice_transition_8665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 558_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3817_branch_ack_1, ack => zeropad3D_CP_2152_elements(558)); -- 
    -- CP-element group 559:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	557 
    -- CP-element group 559: successors 
    -- CP-element group 559: 	560 
    -- CP-element group 559: 	561 
    -- CP-element group 559: 	563 
    -- CP-element group 559:  members (27) 
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842__entry__
      -- CP-element group 559: 	 branch_block_stmt_714/merge_stmt_3823__exit__
      -- CP-element group 559: 	 branch_block_stmt_714/if_stmt_3817_else_link/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/if_stmt_3817_else_link/else_choice_transition
      -- CP-element group 559: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_lorx_xlhsx_xfalse1148
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_sample_start_
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_update_start_
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_word_address_calculated
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_root_address_calculated
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/word_access_start/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/word_access_start/word_0/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/word_access_start/word_0/rr
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/word_access_complete/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/word_access_complete/word_0/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/word_access_complete/word_0/cr
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_update_start_
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Update/cr
      -- CP-element group 559: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_lorx_xlhsx_xfalse1148_PhiReq/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1141_lorx_xlhsx_xfalse1148_PhiReq/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/merge_stmt_3823_PhiReqMerge
      -- CP-element group 559: 	 branch_block_stmt_714/merge_stmt_3823_PhiAck/$entry
      -- CP-element group 559: 	 branch_block_stmt_714/merge_stmt_3823_PhiAck/$exit
      -- CP-element group 559: 	 branch_block_stmt_714/merge_stmt_3823_PhiAck/dummy
      -- 
    else_choice_transition_8669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3817_branch_ack_0, ack => zeropad3D_CP_2152_elements(559)); -- 
    rr_8690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(559), ack => LOAD_col_high_3825_load_0_req_0); -- 
    cr_8701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(559), ack => LOAD_col_high_3825_load_0_req_1); -- 
    cr_8720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(559), ack => type_cast_3829_inst_req_1); -- 
    -- CP-element group 560:  transition  input  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	559 
    -- CP-element group 560: successors 
    -- CP-element group 560:  members (5) 
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_sample_completed_
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/$exit
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/word_access_start/$exit
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/word_access_start/word_0/$exit
      -- CP-element group 560: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Sample/word_access_start/word_0/ra
      -- 
    ra_8691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3825_load_0_ack_0, ack => zeropad3D_CP_2152_elements(560)); -- 
    -- CP-element group 561:  transition  input  output  bypass 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	559 
    -- CP-element group 561: successors 
    -- CP-element group 561: 	562 
    -- CP-element group 561:  members (12) 
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_update_completed_
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/word_access_complete/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/word_access_complete/word_0/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/word_access_complete/word_0/ca
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/LOAD_col_high_3825_Merge/$entry
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/LOAD_col_high_3825_Merge/$exit
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/LOAD_col_high_3825_Merge/merge_req
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/LOAD_col_high_3825_Update/LOAD_col_high_3825_Merge/merge_ack
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_sample_start_
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Sample/$entry
      -- CP-element group 561: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Sample/rr
      -- 
    ca_8702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_3825_load_0_ack_1, ack => zeropad3D_CP_2152_elements(561)); -- 
    rr_8715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(561), ack => type_cast_3829_inst_req_0); -- 
    -- CP-element group 562:  transition  input  bypass 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	561 
    -- CP-element group 562: successors 
    -- CP-element group 562:  members (3) 
      -- CP-element group 562: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_sample_completed_
      -- CP-element group 562: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Sample/$exit
      -- CP-element group 562: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Sample/ra
      -- 
    ra_8716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 562_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3829_inst_ack_0, ack => zeropad3D_CP_2152_elements(562)); -- 
    -- CP-element group 563:  branch  transition  place  input  output  bypass 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	559 
    -- CP-element group 563: successors 
    -- CP-element group 563: 	564 
    -- CP-element group 563: 	565 
    -- CP-element group 563:  members (13) 
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842__exit__
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843__entry__
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/$exit
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_update_completed_
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Update/$exit
      -- CP-element group 563: 	 branch_block_stmt_714/assign_stmt_3826_to_assign_stmt_3842/type_cast_3829_Update/ca
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843_dead_link/$entry
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843_eval_test/$entry
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843_eval_test/$exit
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843_eval_test/branch_req
      -- CP-element group 563: 	 branch_block_stmt_714/R_cmp1156_3844_place
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843_if_link/$entry
      -- CP-element group 563: 	 branch_block_stmt_714/if_stmt_3843_else_link/$entry
      -- 
    ca_8721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 563_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3829_inst_ack_1, ack => zeropad3D_CP_2152_elements(563)); -- 
    branch_req_8729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(563), ack => if_stmt_3843_branch_req_0); -- 
    -- CP-element group 564:  fork  transition  place  input  output  bypass 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	563 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	580 
    -- CP-element group 564: 	581 
    -- CP-element group 564: 	583 
    -- CP-element group 564: 	585 
    -- CP-element group 564: 	587 
    -- CP-element group 564: 	589 
    -- CP-element group 564: 	591 
    -- CP-element group 564: 	593 
    -- CP-element group 564: 	595 
    -- CP-element group 564: 	598 
    -- CP-element group 564:  members (46) 
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012__entry__
      -- CP-element group 564: 	 branch_block_stmt_714/merge_stmt_3907__exit__
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/word_access_complete/word_0/cr
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_update_start
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Update/cr
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_complete/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_complete/req
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Update/req
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/word_access_complete/word_0/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/word_access_complete/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_complete/req
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Update/req
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_update_start
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_complete/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/if_stmt_3843_if_link/$exit
      -- CP-element group 564: 	 branch_block_stmt_714/if_stmt_3843_if_link/if_choice_transition
      -- CP-element group 564: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xelse1179
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_sample_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Sample/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Sample/rr
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Update/cr
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Update/cr
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_update_start_
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/word_access_complete/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/word_access_complete/word_0/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/word_access_complete/word_0/cr
      -- CP-element group 564: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xelse1179_PhiReq/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xelse1179_PhiReq/$exit
      -- CP-element group 564: 	 branch_block_stmt_714/merge_stmt_3907_PhiReqMerge
      -- CP-element group 564: 	 branch_block_stmt_714/merge_stmt_3907_PhiAck/$entry
      -- CP-element group 564: 	 branch_block_stmt_714/merge_stmt_3907_PhiAck/$exit
      -- CP-element group 564: 	 branch_block_stmt_714/merge_stmt_3907_PhiAck/dummy
      -- 
    if_choice_transition_8734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 564_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3843_branch_ack_1, ack => zeropad3D_CP_2152_elements(564)); -- 
    cr_9002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => ptr_deref_3986_load_0_req_1); -- 
    cr_9021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => type_cast_4000_inst_req_1); -- 
    req_8957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => addr_of_3982_final_reg_req_1); -- 
    req_9052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => array_obj_ref_4006_index_offset_req_1); -- 
    req_9067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => addr_of_4007_final_reg_req_1); -- 
    req_8942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => array_obj_ref_3981_index_offset_req_1); -- 
    rr_8892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => type_cast_3911_inst_req_0); -- 
    cr_8897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => type_cast_3911_inst_req_1); -- 
    cr_8911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => type_cast_3975_inst_req_1); -- 
    cr_9117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(564), ack => ptr_deref_4010_store_0_req_1); -- 
    -- CP-element group 565:  transition  place  input  bypass 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	563 
    -- CP-element group 565: successors 
    -- CP-element group 565: 	1073 
    -- CP-element group 565:  members (5) 
      -- CP-element group 565: 	 branch_block_stmt_714/if_stmt_3843_else_link/$exit
      -- CP-element group 565: 	 branch_block_stmt_714/if_stmt_3843_else_link/else_choice_transition
      -- CP-element group 565: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xthen1158
      -- CP-element group 565: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xthen1158_PhiReq/$entry
      -- CP-element group 565: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1148_ifx_xthen1158_PhiReq/$exit
      -- 
    else_choice_transition_8738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3843_branch_ack_0, ack => zeropad3D_CP_2152_elements(565)); -- 
    -- CP-element group 566:  transition  input  bypass 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	1073 
    -- CP-element group 566: successors 
    -- CP-element group 566:  members (3) 
      -- CP-element group 566: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_sample_completed_
      -- CP-element group 566: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Sample/$exit
      -- CP-element group 566: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Sample/ra
      -- 
    ra_8752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 566_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3853_inst_ack_0, ack => zeropad3D_CP_2152_elements(566)); -- 
    -- CP-element group 567:  transition  input  bypass 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	1073 
    -- CP-element group 567: successors 
    -- CP-element group 567: 	570 
    -- CP-element group 567:  members (3) 
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_update_completed_
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Update/$exit
      -- CP-element group 567: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Update/ca
      -- 
    ca_8757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3853_inst_ack_1, ack => zeropad3D_CP_2152_elements(567)); -- 
    -- CP-element group 568:  transition  input  bypass 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	1073 
    -- CP-element group 568: successors 
    -- CP-element group 568:  members (3) 
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_sample_completed_
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Sample/$exit
      -- CP-element group 568: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Sample/ra
      -- 
    ra_8766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 568_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3858_inst_ack_0, ack => zeropad3D_CP_2152_elements(568)); -- 
    -- CP-element group 569:  transition  input  bypass 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	1073 
    -- CP-element group 569: successors 
    -- CP-element group 569: 	570 
    -- CP-element group 569:  members (3) 
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_update_completed_
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Update/$exit
      -- CP-element group 569: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Update/ca
      -- 
    ca_8771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 569_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3858_inst_ack_1, ack => zeropad3D_CP_2152_elements(569)); -- 
    -- CP-element group 570:  join  transition  output  bypass 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	567 
    -- CP-element group 570: 	569 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	571 
    -- CP-element group 570:  members (3) 
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_sample_start_
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Sample/$entry
      -- CP-element group 570: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Sample/rr
      -- 
    rr_8779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(570), ack => type_cast_3892_inst_req_0); -- 
    zeropad3D_cp_element_group_570: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_570"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(567) & zeropad3D_CP_2152_elements(569);
      gj_zeropad3D_cp_element_group_570 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(570), clk => clk, reset => reset); --
    end block;
    -- CP-element group 571:  transition  input  bypass 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	570 
    -- CP-element group 571: successors 
    -- CP-element group 571:  members (3) 
      -- CP-element group 571: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_sample_completed_
      -- CP-element group 571: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Sample/$exit
      -- CP-element group 571: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Sample/ra
      -- 
    ra_8780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 571_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3892_inst_ack_0, ack => zeropad3D_CP_2152_elements(571)); -- 
    -- CP-element group 572:  transition  input  output  bypass 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	1073 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	573 
    -- CP-element group 572:  members (16) 
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_update_completed_
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Update/$exit
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Update/ca
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_resized_1
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_scaled_1
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_computed_1
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_resize_1/$entry
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_resize_1/$exit
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_resize_1/index_resize_req
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_resize_1/index_resize_ack
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_scale_1/$entry
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_scale_1/$exit
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_scale_1/scale_rename_req
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_index_scale_1/scale_rename_ack
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Sample/$entry
      -- CP-element group 572: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Sample/req
      -- 
    ca_8785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3892_inst_ack_1, ack => zeropad3D_CP_2152_elements(572)); -- 
    req_8810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(572), ack => array_obj_ref_3898_index_offset_req_0); -- 
    -- CP-element group 573:  transition  input  bypass 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	572 
    -- CP-element group 573: successors 
    -- CP-element group 573: 	579 
    -- CP-element group 573:  members (3) 
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_sample_complete
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Sample/$exit
      -- CP-element group 573: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Sample/ack
      -- 
    ack_8811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 573_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3898_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(573)); -- 
    -- CP-element group 574:  transition  input  output  bypass 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	1073 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	575 
    -- CP-element group 574:  members (11) 
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_sample_start_
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_root_address_calculated
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_offset_calculated
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Update/$exit
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Update/ack
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_base_plus_offset/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_base_plus_offset/$exit
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_base_plus_offset/sum_rename_req
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_base_plus_offset/sum_rename_ack
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_request/$entry
      -- CP-element group 574: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_request/req
      -- 
    ack_8816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3898_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(574)); -- 
    req_8825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(574), ack => addr_of_3899_final_reg_req_0); -- 
    -- CP-element group 575:  transition  input  bypass 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	574 
    -- CP-element group 575: successors 
    -- CP-element group 575:  members (3) 
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_sample_completed_
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_request/$exit
      -- CP-element group 575: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_request/ack
      -- 
    ack_8826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3899_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(575)); -- 
    -- CP-element group 576:  join  fork  transition  input  output  bypass 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	1073 
    -- CP-element group 576: successors 
    -- CP-element group 576: 	577 
    -- CP-element group 576:  members (28) 
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_update_completed_
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_complete/$exit
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_complete/ack
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_sample_start_
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_address_calculated
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_word_address_calculated
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_root_address_calculated
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_address_resized
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_addr_resize/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_addr_resize/$exit
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_addr_resize/base_resize_req
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_addr_resize/base_resize_ack
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_plus_offset/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_plus_offset/$exit
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_plus_offset/sum_rename_req
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_base_plus_offset/sum_rename_ack
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_word_addrgen/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_word_addrgen/$exit
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_word_addrgen/root_register_req
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_word_addrgen/root_register_ack
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/ptr_deref_3902_Split/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/ptr_deref_3902_Split/$exit
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/ptr_deref_3902_Split/split_req
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/ptr_deref_3902_Split/split_ack
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/word_access_start/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/word_access_start/word_0/$entry
      -- CP-element group 576: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/word_access_start/word_0/rr
      -- 
    ack_8831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3899_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(576)); -- 
    rr_8869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(576), ack => ptr_deref_3902_store_0_req_0); -- 
    -- CP-element group 577:  transition  input  bypass 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	576 
    -- CP-element group 577: successors 
    -- CP-element group 577:  members (5) 
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_sample_completed_
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/$exit
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/word_access_start/$exit
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/word_access_start/word_0/$exit
      -- CP-element group 577: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Sample/word_access_start/word_0/ra
      -- 
    ra_8870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 577_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3902_store_0_ack_0, ack => zeropad3D_CP_2152_elements(577)); -- 
    -- CP-element group 578:  transition  input  bypass 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	1073 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	579 
    -- CP-element group 578:  members (5) 
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_update_completed_
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/$exit
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/word_access_complete/$exit
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/word_access_complete/word_0/$exit
      -- CP-element group 578: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/word_access_complete/word_0/ca
      -- 
    ca_8881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 578_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3902_store_0_ack_1, ack => zeropad3D_CP_2152_elements(578)); -- 
    -- CP-element group 579:  join  transition  place  bypass 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	573 
    -- CP-element group 579: 	578 
    -- CP-element group 579: successors 
    -- CP-element group 579: 	1074 
    -- CP-element group 579:  members (5) 
      -- CP-element group 579: 	 branch_block_stmt_714/ifx_xthen1158_ifx_xend1227
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905__exit__
      -- CP-element group 579: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/$exit
      -- CP-element group 579: 	 branch_block_stmt_714/ifx_xthen1158_ifx_xend1227_PhiReq/$entry
      -- CP-element group 579: 	 branch_block_stmt_714/ifx_xthen1158_ifx_xend1227_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_579: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_579"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(573) & zeropad3D_CP_2152_elements(578);
      gj_zeropad3D_cp_element_group_579 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(579), clk => clk, reset => reset); --
    end block;
    -- CP-element group 580:  transition  input  bypass 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	564 
    -- CP-element group 580: successors 
    -- CP-element group 580:  members (3) 
      -- CP-element group 580: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_sample_completed_
      -- CP-element group 580: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Sample/$exit
      -- CP-element group 580: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Sample/ra
      -- 
    ra_8893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3911_inst_ack_0, ack => zeropad3D_CP_2152_elements(580)); -- 
    -- CP-element group 581:  fork  transition  input  output  bypass 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	564 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	582 
    -- CP-element group 581: 	590 
    -- CP-element group 581:  members (9) 
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_sample_start_
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Sample/$entry
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Sample/rr
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_update_completed_
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Update/$exit
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3911_Update/ca
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_sample_start_
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Sample/$entry
      -- CP-element group 581: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Sample/rr
      -- 
    ca_8898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 581_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3911_inst_ack_1, ack => zeropad3D_CP_2152_elements(581)); -- 
    rr_8906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(581), ack => type_cast_3975_inst_req_0); -- 
    rr_9016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(581), ack => type_cast_4000_inst_req_0); -- 
    -- CP-element group 582:  transition  input  bypass 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	581 
    -- CP-element group 582: successors 
    -- CP-element group 582:  members (3) 
      -- CP-element group 582: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_sample_completed_
      -- CP-element group 582: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Sample/$exit
      -- CP-element group 582: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Sample/ra
      -- 
    ra_8907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 582_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3975_inst_ack_0, ack => zeropad3D_CP_2152_elements(582)); -- 
    -- CP-element group 583:  transition  input  output  bypass 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	564 
    -- CP-element group 583: successors 
    -- CP-element group 583: 	584 
    -- CP-element group 583:  members (16) 
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_resized_1
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_scaled_1
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_computed_1
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_resize_1/$entry
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_resize_1/$exit
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_resize_1/index_resize_req
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_resize_1/index_resize_ack
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_scale_1/$entry
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_scale_1/$exit
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Sample/req
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Sample/$entry
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_scale_1/scale_rename_ack
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_index_scale_1/scale_rename_req
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_update_completed_
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Update/$exit
      -- CP-element group 583: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_3975_Update/ca
      -- 
    ca_8912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3975_inst_ack_1, ack => zeropad3D_CP_2152_elements(583)); -- 
    req_8937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(583), ack => array_obj_ref_3981_index_offset_req_0); -- 
    -- CP-element group 584:  transition  input  bypass 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	583 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	599 
    -- CP-element group 584:  members (3) 
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Sample/ack
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Sample/$exit
      -- CP-element group 584: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_sample_complete
      -- 
    ack_8938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 584_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3981_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(584)); -- 
    -- CP-element group 585:  transition  input  output  bypass 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	564 
    -- CP-element group 585: successors 
    -- CP-element group 585: 	586 
    -- CP-element group 585:  members (11) 
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_base_plus_offset/$entry
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_base_plus_offset/$exit
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_base_plus_offset/sum_rename_req
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_base_plus_offset/sum_rename_ack
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_request/$entry
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_offset_calculated
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Update/ack
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_final_index_sum_regn_Update/$exit
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_3981_root_address_calculated
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_request/req
      -- CP-element group 585: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_sample_start_
      -- 
    ack_8943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 585_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3981_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(585)); -- 
    req_8952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(585), ack => addr_of_3982_final_reg_req_0); -- 
    -- CP-element group 586:  transition  input  bypass 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	585 
    -- CP-element group 586: successors 
    -- CP-element group 586:  members (3) 
      -- CP-element group 586: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_request/ack
      -- CP-element group 586: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_request/$exit
      -- CP-element group 586: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_sample_completed_
      -- 
    ack_8953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 586_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3982_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(586)); -- 
    -- CP-element group 587:  join  fork  transition  input  output  bypass 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	564 
    -- CP-element group 587: successors 
    -- CP-element group 587: 	588 
    -- CP-element group 587:  members (24) 
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_complete/$exit
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_root_address_calculated
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_complete/ack
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_address_resized
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_sample_start_
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_addr_resize/$entry
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/word_access_start/word_0/rr
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/word_access_start/word_0/$entry
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/word_access_start/$entry
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/$entry
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_word_addrgen/root_register_ack
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_word_addrgen/root_register_req
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_word_address_calculated
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_word_addrgen/$exit
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_3982_update_completed_
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_address_calculated
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_word_addrgen/$entry
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_plus_offset/sum_rename_ack
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_plus_offset/sum_rename_req
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_plus_offset/$exit
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_plus_offset/$entry
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_addr_resize/base_resize_ack
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_addr_resize/base_resize_req
      -- CP-element group 587: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_base_addr_resize/$exit
      -- 
    ack_8958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 587_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3982_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(587)); -- 
    rr_8991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(587), ack => ptr_deref_3986_load_0_req_0); -- 
    -- CP-element group 588:  transition  input  bypass 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	587 
    -- CP-element group 588: successors 
    -- CP-element group 588:  members (5) 
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_sample_completed_
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/word_access_start/word_0/ra
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/word_access_start/word_0/$exit
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/word_access_start/$exit
      -- CP-element group 588: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Sample/$exit
      -- 
    ra_8992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3986_load_0_ack_0, ack => zeropad3D_CP_2152_elements(588)); -- 
    -- CP-element group 589:  transition  input  bypass 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	564 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	596 
    -- CP-element group 589:  members (9) 
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/word_access_complete/word_0/$exit
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/word_access_complete/word_0/ca
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/ptr_deref_3986_Merge/$entry
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/ptr_deref_3986_Merge/$exit
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/ptr_deref_3986_Merge/merge_req
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/ptr_deref_3986_Merge/merge_ack
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/word_access_complete/$exit
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_Update/$exit
      -- CP-element group 589: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_3986_update_completed_
      -- 
    ca_9003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 589_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3986_load_0_ack_1, ack => zeropad3D_CP_2152_elements(589)); -- 
    -- CP-element group 590:  transition  input  bypass 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	581 
    -- CP-element group 590: successors 
    -- CP-element group 590:  members (3) 
      -- CP-element group 590: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_sample_completed_
      -- CP-element group 590: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Sample/$exit
      -- CP-element group 590: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Sample/ra
      -- 
    ra_9017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 590_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4000_inst_ack_0, ack => zeropad3D_CP_2152_elements(590)); -- 
    -- CP-element group 591:  transition  input  output  bypass 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	564 
    -- CP-element group 591: successors 
    -- CP-element group 591: 	592 
    -- CP-element group 591:  members (16) 
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Sample/$entry
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Update/ca
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Sample/req
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_update_completed_
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_resized_1
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/type_cast_4000_Update/$exit
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_scale_1/scale_rename_ack
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_scale_1/scale_rename_req
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_scale_1/$exit
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_scale_1/$entry
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_resize_1/index_resize_ack
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_resize_1/index_resize_req
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_resize_1/$exit
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_resize_1/$entry
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_computed_1
      -- CP-element group 591: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_index_scaled_1
      -- 
    ca_9022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 591_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4000_inst_ack_1, ack => zeropad3D_CP_2152_elements(591)); -- 
    req_9047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(591), ack => array_obj_ref_4006_index_offset_req_0); -- 
    -- CP-element group 592:  transition  input  bypass 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	591 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	599 
    -- CP-element group 592:  members (3) 
      -- CP-element group 592: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Sample/$exit
      -- CP-element group 592: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Sample/ack
      -- CP-element group 592: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_sample_complete
      -- 
    ack_9048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4006_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(592)); -- 
    -- CP-element group 593:  transition  input  output  bypass 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	564 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	594 
    -- CP-element group 593:  members (11) 
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_request/$entry
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_request/req
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_sample_start_
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Update/$exit
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_root_address_calculated
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_offset_calculated
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_final_index_sum_regn_Update/ack
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_base_plus_offset/sum_rename_ack
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_base_plus_offset/sum_rename_req
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_base_plus_offset/$exit
      -- CP-element group 593: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/array_obj_ref_4006_base_plus_offset/$entry
      -- 
    ack_9053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 593_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4006_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(593)); -- 
    req_9062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(593), ack => addr_of_4007_final_reg_req_0); -- 
    -- CP-element group 594:  transition  input  bypass 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	593 
    -- CP-element group 594: successors 
    -- CP-element group 594:  members (3) 
      -- CP-element group 594: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_request/$exit
      -- CP-element group 594: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_request/ack
      -- CP-element group 594: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_sample_completed_
      -- 
    ack_9063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 594_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4007_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(594)); -- 
    -- CP-element group 595:  fork  transition  input  bypass 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	564 
    -- CP-element group 595: successors 
    -- CP-element group 595: 	596 
    -- CP-element group 595:  members (19) 
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_complete/ack
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_word_addrgen/root_register_req
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_addr_resize/base_resize_req
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_word_address_calculated
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_addr_resize/base_resize_ack
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_plus_offset/$entry
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_word_addrgen/root_register_ack
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_plus_offset/$exit
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_complete/$exit
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/addr_of_4007_update_completed_
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_address_calculated
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_word_addrgen/$exit
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_word_addrgen/$entry
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_plus_offset/sum_rename_ack
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_addr_resize/$exit
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_plus_offset/sum_rename_req
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_addr_resize/$entry
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_base_address_resized
      -- CP-element group 595: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_root_address_calculated
      -- 
    ack_9068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4007_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(595)); -- 
    -- CP-element group 596:  join  transition  output  bypass 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	589 
    -- CP-element group 596: 	595 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	597 
    -- CP-element group 596:  members (9) 
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_sample_start_
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/ptr_deref_4010_Split/$entry
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/ptr_deref_4010_Split/$exit
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/$entry
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/ptr_deref_4010_Split/split_req
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/ptr_deref_4010_Split/split_ack
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/word_access_start/$entry
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/word_access_start/word_0/$entry
      -- CP-element group 596: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/word_access_start/word_0/rr
      -- 
    rr_9106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(596), ack => ptr_deref_4010_store_0_req_0); -- 
    zeropad3D_cp_element_group_596: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_596"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(589) & zeropad3D_CP_2152_elements(595);
      gj_zeropad3D_cp_element_group_596 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(596), clk => clk, reset => reset); --
    end block;
    -- CP-element group 597:  transition  input  bypass 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	596 
    -- CP-element group 597: successors 
    -- CP-element group 597:  members (5) 
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_sample_completed_
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/word_access_start/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/word_access_start/word_0/$exit
      -- CP-element group 597: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Sample/word_access_start/word_0/ra
      -- 
    ra_9107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 597_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4010_store_0_ack_0, ack => zeropad3D_CP_2152_elements(597)); -- 
    -- CP-element group 598:  transition  input  bypass 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	564 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	599 
    -- CP-element group 598:  members (5) 
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_update_completed_
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/$exit
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/word_access_complete/$exit
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/word_access_complete/word_0/$exit
      -- CP-element group 598: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/ptr_deref_4010_Update/word_access_complete/word_0/ca
      -- 
    ca_9118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 598_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4010_store_0_ack_1, ack => zeropad3D_CP_2152_elements(598)); -- 
    -- CP-element group 599:  join  transition  place  bypass 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	584 
    -- CP-element group 599: 	592 
    -- CP-element group 599: 	598 
    -- CP-element group 599: successors 
    -- CP-element group 599: 	1074 
    -- CP-element group 599:  members (5) 
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012__exit__
      -- CP-element group 599: 	 branch_block_stmt_714/ifx_xelse1179_ifx_xend1227
      -- CP-element group 599: 	 branch_block_stmt_714/assign_stmt_3912_to_assign_stmt_4012/$exit
      -- CP-element group 599: 	 branch_block_stmt_714/ifx_xelse1179_ifx_xend1227_PhiReq/$entry
      -- CP-element group 599: 	 branch_block_stmt_714/ifx_xelse1179_ifx_xend1227_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_599: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_599"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(584) & zeropad3D_CP_2152_elements(592) & zeropad3D_CP_2152_elements(598);
      gj_zeropad3D_cp_element_group_599 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(599), clk => clk, reset => reset); --
    end block;
    -- CP-element group 600:  transition  input  bypass 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	1074 
    -- CP-element group 600: successors 
    -- CP-element group 600:  members (3) 
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_sample_completed_
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Sample/$exit
      -- CP-element group 600: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Sample/ra
      -- 
    ra_9130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4018_inst_ack_0, ack => zeropad3D_CP_2152_elements(600)); -- 
    -- CP-element group 601:  branch  transition  place  input  output  bypass 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	1074 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	602 
    -- CP-element group 601: 	603 
    -- CP-element group 601:  members (13) 
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032__exit__
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033__entry__
      -- CP-element group 601: 	 branch_block_stmt_714/R_cmp1235_4034_place
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_update_completed_
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Update/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Update/ca
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033_dead_link/$entry
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033_eval_test/$entry
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033_eval_test/$exit
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033_eval_test/branch_req
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033_if_link/$entry
      -- CP-element group 601: 	 branch_block_stmt_714/if_stmt_4033_else_link/$entry
      -- 
    ca_9135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 601_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4018_inst_ack_1, ack => zeropad3D_CP_2152_elements(601)); -- 
    branch_req_9143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(601), ack => if_stmt_4033_branch_req_0); -- 
    -- CP-element group 602:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	601 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	1083 
    -- CP-element group 602: 	1084 
    -- CP-element group 602: 	1086 
    -- CP-element group 602: 	1087 
    -- CP-element group 602: 	1089 
    -- CP-element group 602: 	1090 
    -- CP-element group 602:  members (40) 
      -- CP-element group 602: 	 branch_block_stmt_714/merge_stmt_4039__exit__
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4045__entry__
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4045__exit__
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xend1227_ifx_xthen1237
      -- CP-element group 602: 	 branch_block_stmt_714/if_stmt_4033_if_link/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/if_stmt_4033_if_link/if_choice_transition
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4045/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/assign_stmt_4045/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Update/cr
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Update/cr
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Update/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Sample/rr
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Update/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Sample/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Sample/rr
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xend1227_ifx_xthen1237_PhiReq/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xend1227_ifx_xthen1237_PhiReq/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/merge_stmt_4039_PhiReqMerge
      -- CP-element group 602: 	 branch_block_stmt_714/merge_stmt_4039_PhiAck/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/merge_stmt_4039_PhiAck/$exit
      -- CP-element group 602: 	 branch_block_stmt_714/merge_stmt_4039_PhiAck/dummy
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Sample/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Sample/rr
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Update/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Update/cr
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/$entry
      -- CP-element group 602: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Sample/$entry
      -- 
    if_choice_transition_9148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 602_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4033_branch_ack_1, ack => zeropad3D_CP_2152_elements(602)); -- 
    cr_13663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(602), ack => type_cast_4142_inst_req_1); -- 
    cr_13686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(602), ack => type_cast_4148_inst_req_1); -- 
    rr_13681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(602), ack => type_cast_4148_inst_req_0); -- 
    rr_13658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(602), ack => type_cast_4142_inst_req_0); -- 
    rr_13635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(602), ack => type_cast_4135_inst_req_0); -- 
    cr_13640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(602), ack => type_cast_4135_inst_req_1); -- 
    -- CP-element group 603:  fork  transition  place  input  output  bypass 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	601 
    -- CP-element group 603: successors 
    -- CP-element group 603: 	604 
    -- CP-element group 603: 	605 
    -- CP-element group 603: 	606 
    -- CP-element group 603: 	607 
    -- CP-element group 603: 	609 
    -- CP-element group 603: 	612 
    -- CP-element group 603: 	614 
    -- CP-element group 603: 	615 
    -- CP-element group 603: 	616 
    -- CP-element group 603: 	618 
    -- CP-element group 603:  members (54) 
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124__entry__
      -- CP-element group 603: 	 branch_block_stmt_714/merge_stmt_4047__exit__
      -- CP-element group 603: 	 branch_block_stmt_714/ifx_xend1227_ifx_xelse1242
      -- CP-element group 603: 	 branch_block_stmt_714/if_stmt_4033_else_link/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/if_stmt_4033_else_link/else_choice_transition
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_sample_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Sample/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Sample/rr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Update/cr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_sample_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_word_address_calculated
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_root_address_calculated
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/word_access_start/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/word_access_start/word_0/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/word_access_start/word_0/rr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/word_access_complete/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/word_access_complete/word_0/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/word_access_complete/word_0/cr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Update/cr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Update/cr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Update/cr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_sample_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_word_address_calculated
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_root_address_calculated
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/word_access_start/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/word_access_start/word_0/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/word_access_start/word_0/rr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/word_access_complete/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/word_access_complete/word_0/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/word_access_complete/word_0/cr
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_update_start_
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Update/cr
      -- CP-element group 603: 	 branch_block_stmt_714/ifx_xend1227_ifx_xelse1242_PhiReq/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/ifx_xend1227_ifx_xelse1242_PhiReq/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/merge_stmt_4047_PhiReqMerge
      -- CP-element group 603: 	 branch_block_stmt_714/merge_stmt_4047_PhiAck/$entry
      -- CP-element group 603: 	 branch_block_stmt_714/merge_stmt_4047_PhiAck/$exit
      -- CP-element group 603: 	 branch_block_stmt_714/merge_stmt_4047_PhiAck/dummy
      -- 
    else_choice_transition_9152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 603_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4033_branch_ack_0, ack => zeropad3D_CP_2152_elements(603)); -- 
    rr_9168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => type_cast_4057_inst_req_0); -- 
    cr_9173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => type_cast_4057_inst_req_1); -- 
    rr_9190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => LOAD_col_high_4060_load_0_req_0); -- 
    cr_9201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => LOAD_col_high_4060_load_0_req_1); -- 
    cr_9220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => type_cast_4064_inst_req_1); -- 
    cr_9234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => type_cast_4078_inst_req_1); -- 
    cr_9248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => type_cast_4094_inst_req_1); -- 
    rr_9265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => LOAD_row_high_4097_load_0_req_0); -- 
    cr_9276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => LOAD_row_high_4097_load_0_req_1); -- 
    cr_9295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(603), ack => type_cast_4101_inst_req_1); -- 
    -- CP-element group 604:  transition  input  bypass 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	603 
    -- CP-element group 604: successors 
    -- CP-element group 604:  members (3) 
      -- CP-element group 604: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_sample_completed_
      -- CP-element group 604: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Sample/$exit
      -- CP-element group 604: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Sample/ra
      -- 
    ra_9169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 604_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4057_inst_ack_0, ack => zeropad3D_CP_2152_elements(604)); -- 
    -- CP-element group 605:  transition  input  bypass 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	603 
    -- CP-element group 605: successors 
    -- CP-element group 605: 	610 
    -- CP-element group 605:  members (3) 
      -- CP-element group 605: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_update_completed_
      -- CP-element group 605: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Update/$exit
      -- CP-element group 605: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4057_Update/ca
      -- 
    ca_9174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 605_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4057_inst_ack_1, ack => zeropad3D_CP_2152_elements(605)); -- 
    -- CP-element group 606:  transition  input  bypass 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	603 
    -- CP-element group 606: successors 
    -- CP-element group 606:  members (5) 
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_sample_completed_
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/$exit
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/word_access_start/$exit
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/word_access_start/word_0/$exit
      -- CP-element group 606: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Sample/word_access_start/word_0/ra
      -- 
    ra_9191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 606_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4060_load_0_ack_0, ack => zeropad3D_CP_2152_elements(606)); -- 
    -- CP-element group 607:  transition  input  output  bypass 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	603 
    -- CP-element group 607: successors 
    -- CP-element group 607: 	608 
    -- CP-element group 607:  members (12) 
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_update_completed_
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/$exit
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/word_access_complete/$exit
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/word_access_complete/word_0/$exit
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/word_access_complete/word_0/ca
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/LOAD_col_high_4060_Merge/$entry
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/LOAD_col_high_4060_Merge/$exit
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/LOAD_col_high_4060_Merge/merge_req
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_col_high_4060_Update/LOAD_col_high_4060_Merge/merge_ack
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_sample_start_
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Sample/$entry
      -- CP-element group 607: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Sample/rr
      -- 
    ca_9202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4060_load_0_ack_1, ack => zeropad3D_CP_2152_elements(607)); -- 
    rr_9215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(607), ack => type_cast_4064_inst_req_0); -- 
    -- CP-element group 608:  transition  input  bypass 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	607 
    -- CP-element group 608: successors 
    -- CP-element group 608:  members (3) 
      -- CP-element group 608: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_sample_completed_
      -- CP-element group 608: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Sample/$exit
      -- CP-element group 608: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Sample/ra
      -- 
    ra_9216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 608_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4064_inst_ack_0, ack => zeropad3D_CP_2152_elements(608)); -- 
    -- CP-element group 609:  transition  input  bypass 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	603 
    -- CP-element group 609: successors 
    -- CP-element group 609: 	610 
    -- CP-element group 609:  members (3) 
      -- CP-element group 609: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_update_completed_
      -- CP-element group 609: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Update/$exit
      -- CP-element group 609: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4064_Update/ca
      -- 
    ca_9221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 609_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4064_inst_ack_1, ack => zeropad3D_CP_2152_elements(609)); -- 
    -- CP-element group 610:  join  transition  output  bypass 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	605 
    -- CP-element group 610: 	609 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	611 
    -- CP-element group 610:  members (3) 
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_sample_start_
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Sample/$entry
      -- CP-element group 610: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Sample/rr
      -- 
    rr_9229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(610), ack => type_cast_4078_inst_req_0); -- 
    zeropad3D_cp_element_group_610: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_610"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(605) & zeropad3D_CP_2152_elements(609);
      gj_zeropad3D_cp_element_group_610 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(610), clk => clk, reset => reset); --
    end block;
    -- CP-element group 611:  transition  input  bypass 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	610 
    -- CP-element group 611: successors 
    -- CP-element group 611:  members (3) 
      -- CP-element group 611: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_sample_completed_
      -- CP-element group 611: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Sample/$exit
      -- CP-element group 611: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Sample/ra
      -- 
    ra_9230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 611_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4078_inst_ack_0, ack => zeropad3D_CP_2152_elements(611)); -- 
    -- CP-element group 612:  transition  input  output  bypass 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	603 
    -- CP-element group 612: successors 
    -- CP-element group 612: 	613 
    -- CP-element group 612:  members (6) 
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_update_completed_
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Update/$exit
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4078_Update/ca
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_sample_start_
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Sample/$entry
      -- CP-element group 612: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Sample/rr
      -- 
    ca_9235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 612_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4078_inst_ack_1, ack => zeropad3D_CP_2152_elements(612)); -- 
    rr_9243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(612), ack => type_cast_4094_inst_req_0); -- 
    -- CP-element group 613:  transition  input  bypass 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	612 
    -- CP-element group 613: successors 
    -- CP-element group 613:  members (3) 
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_sample_completed_
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Sample/$exit
      -- CP-element group 613: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Sample/ra
      -- 
    ra_9244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 613_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4094_inst_ack_0, ack => zeropad3D_CP_2152_elements(613)); -- 
    -- CP-element group 614:  transition  input  bypass 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	603 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	619 
    -- CP-element group 614:  members (3) 
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_update_completed_
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Update/$exit
      -- CP-element group 614: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4094_Update/ca
      -- 
    ca_9249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 614_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4094_inst_ack_1, ack => zeropad3D_CP_2152_elements(614)); -- 
    -- CP-element group 615:  transition  input  bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	603 
    -- CP-element group 615: successors 
    -- CP-element group 615:  members (5) 
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_sample_completed_
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/$exit
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/word_access_start/$exit
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/word_access_start/word_0/$exit
      -- CP-element group 615: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Sample/word_access_start/word_0/ra
      -- 
    ra_9266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4097_load_0_ack_0, ack => zeropad3D_CP_2152_elements(615)); -- 
    -- CP-element group 616:  transition  input  output  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	603 
    -- CP-element group 616: successors 
    -- CP-element group 616: 	617 
    -- CP-element group 616:  members (12) 
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_update_completed_
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/word_access_complete/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/word_access_complete/word_0/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/word_access_complete/word_0/ca
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/LOAD_row_high_4097_Merge/$entry
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/LOAD_row_high_4097_Merge/$exit
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/LOAD_row_high_4097_Merge/merge_req
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/LOAD_row_high_4097_Update/LOAD_row_high_4097_Merge/merge_ack
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_sample_start_
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Sample/$entry
      -- CP-element group 616: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Sample/rr
      -- 
    ca_9277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 616_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4097_load_0_ack_1, ack => zeropad3D_CP_2152_elements(616)); -- 
    rr_9290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(616), ack => type_cast_4101_inst_req_0); -- 
    -- CP-element group 617:  transition  input  bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	616 
    -- CP-element group 617: successors 
    -- CP-element group 617:  members (3) 
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_sample_completed_
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Sample/$exit
      -- CP-element group 617: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Sample/ra
      -- 
    ra_9291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4101_inst_ack_0, ack => zeropad3D_CP_2152_elements(617)); -- 
    -- CP-element group 618:  transition  input  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	603 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	619 
    -- CP-element group 618:  members (3) 
      -- CP-element group 618: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_update_completed_
      -- CP-element group 618: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Update/$exit
      -- CP-element group 618: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/type_cast_4101_Update/ca
      -- 
    ca_9296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 618_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4101_inst_ack_1, ack => zeropad3D_CP_2152_elements(618)); -- 
    -- CP-element group 619:  branch  join  transition  place  output  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	614 
    -- CP-element group 619: 	618 
    -- CP-element group 619: successors 
    -- CP-element group 619: 	620 
    -- CP-element group 619: 	621 
    -- CP-element group 619:  members (10) 
      -- CP-element group 619: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124__exit__
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125__entry__
      -- CP-element group 619: 	 branch_block_stmt_714/R_cmp1270_4126_place
      -- CP-element group 619: 	 branch_block_stmt_714/assign_stmt_4053_to_assign_stmt_4124/$exit
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125_dead_link/$entry
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125_eval_test/$entry
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125_eval_test/$exit
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125_eval_test/branch_req
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125_if_link/$entry
      -- CP-element group 619: 	 branch_block_stmt_714/if_stmt_4125_else_link/$entry
      -- 
    branch_req_9304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(619), ack => if_stmt_4125_branch_req_0); -- 
    zeropad3D_cp_element_group_619: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_619"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(614) & zeropad3D_CP_2152_elements(618);
      gj_zeropad3D_cp_element_group_619 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(619), clk => clk, reset => reset); --
    end block;
    -- CP-element group 620:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	619 
    -- CP-element group 620: successors 
    -- CP-element group 620: 	622 
    -- CP-element group 620: 	623 
    -- CP-element group 620: 	625 
    -- CP-element group 620: 	626 
    -- CP-element group 620: 	627 
    -- CP-element group 620: 	628 
    -- CP-element group 620: 	629 
    -- CP-element group 620: 	630 
    -- CP-element group 620: 	631 
    -- CP-element group 620: 	632 
    -- CP-element group 620: 	633 
    -- CP-element group 620: 	634 
    -- CP-element group 620: 	635 
    -- CP-element group 620: 	637 
    -- CP-element group 620: 	639 
    -- CP-element group 620: 	641 
    -- CP-element group 620:  members (124) 
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294__entry__
      -- CP-element group 620: 	 branch_block_stmt_714/merge_stmt_4153__exit__
      -- CP-element group 620: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4125_if_link/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/if_stmt_4125_if_link/if_choice_transition
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/word_access_complete/word_0/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Update/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/word_access_complete/word_0/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/word_access_complete/word_0/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/word_access_complete/word_0/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_address_resized
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_addr_resize/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_addr_resize/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_addr_resize/base_resize_req
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_addr_resize/base_resize_ack
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_plus_offset/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_plus_offset/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_plus_offset/sum_rename_req
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_base_plus_offset/sum_rename_ack
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_word_addrgen/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_word_addrgen/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_word_addrgen/root_register_req
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_word_addrgen/root_register_ack
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/word_access_complete/word_0/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_word_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_root_address_calculated
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_address_resized
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_addr_resize/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_addr_resize/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_addr_resize/base_resize_req
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_addr_resize/base_resize_ack
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_plus_offset/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_plus_offset/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_plus_offset/sum_rename_req
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_base_plus_offset/sum_rename_ack
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_word_addrgen/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_word_addrgen/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_word_addrgen/root_register_req
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_word_addrgen/root_register_ack
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/word_access_start/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/word_access_start/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/word_access_start/word_0/rr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/word_access_complete/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/word_access_complete/word_0/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/word_access_complete/word_0/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Update/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Update/cr
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_update_start_
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Update/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Update/cr
      -- CP-element group 620: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/merge_stmt_4153_PhiReqMerge
      -- CP-element group 620: 	 branch_block_stmt_714/ifx_xelse1242_whilex_xend1280_PhiReq/$exit
      -- CP-element group 620: 	 branch_block_stmt_714/merge_stmt_4153_PhiAck/$entry
      -- CP-element group 620: 	 branch_block_stmt_714/merge_stmt_4153_PhiAck/dummy
      -- CP-element group 620: 	 branch_block_stmt_714/merge_stmt_4153_PhiAck/$exit
      -- 
    if_choice_transition_9309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4125_branch_ack_1, ack => zeropad3D_CP_2152_elements(620)); -- 
    rr_9334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_row_high_4156_load_0_req_0); -- 
    cr_9345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_row_high_4156_load_0_req_1); -- 
    cr_9364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => type_cast_4160_inst_req_1); -- 
    rr_9381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_pad_4175_load_0_req_0); -- 
    cr_9392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_pad_4175_load_0_req_1); -- 
    rr_9414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_depth_high_4178_load_0_req_0); -- 
    cr_9425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_depth_high_4178_load_0_req_1); -- 
    rr_9447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_col_high_4181_load_0_req_0); -- 
    cr_9458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => LOAD_col_high_4181_load_0_req_1); -- 
    rr_9497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => ptr_deref_4193_load_0_req_0); -- 
    cr_9508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => ptr_deref_4193_load_0_req_1); -- 
    rr_9547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => ptr_deref_4205_load_0_req_0); -- 
    cr_9558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => ptr_deref_4205_load_0_req_1); -- 
    cr_9577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => type_cast_4209_inst_req_1); -- 
    cr_9591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => type_cast_4213_inst_req_1); -- 
    cr_9605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(620), ack => type_cast_4252_inst_req_1); -- 
    -- CP-element group 621:  fork  transition  place  input  output  bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	619 
    -- CP-element group 621: successors 
    -- CP-element group 621: 	1075 
    -- CP-element group 621: 	1076 
    -- CP-element group 621: 	1077 
    -- CP-element group 621: 	1079 
    -- CP-element group 621: 	1080 
    -- CP-element group 621:  members (22) 
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279
      -- CP-element group 621: 	 branch_block_stmt_714/if_stmt_4125_else_link/$exit
      -- CP-element group 621: 	 branch_block_stmt_714/if_stmt_4125_else_link/else_choice_transition
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4132/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Sample/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Sample/rr
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Update/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Update/cr
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Sample/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Sample/rr
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Update/$entry
      -- CP-element group 621: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Update/cr
      -- 
    else_choice_transition_9313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4125_branch_ack_0, ack => zeropad3D_CP_2152_elements(621)); -- 
    rr_13586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(621), ack => type_cast_4144_inst_req_0); -- 
    cr_13591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(621), ack => type_cast_4144_inst_req_1); -- 
    rr_13609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(621), ack => type_cast_4150_inst_req_0); -- 
    cr_13614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(621), ack => type_cast_4150_inst_req_1); -- 
    -- CP-element group 622:  transition  input  bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	620 
    -- CP-element group 622: successors 
    -- CP-element group 622:  members (5) 
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_sample_completed_
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/$exit
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/word_access_start/$exit
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/word_access_start/word_0/$exit
      -- CP-element group 622: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Sample/word_access_start/word_0/ra
      -- 
    ra_9335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 622_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4156_load_0_ack_0, ack => zeropad3D_CP_2152_elements(622)); -- 
    -- CP-element group 623:  transition  input  output  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	620 
    -- CP-element group 623: successors 
    -- CP-element group 623: 	624 
    -- CP-element group 623:  members (12) 
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_update_completed_
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/word_access_complete/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/word_access_complete/word_0/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/word_access_complete/word_0/ca
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/LOAD_row_high_4156_Merge/$entry
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/LOAD_row_high_4156_Merge/$exit
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/LOAD_row_high_4156_Merge/merge_req
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_row_high_4156_Update/LOAD_row_high_4156_Merge/merge_ack
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_sample_start_
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Sample/$entry
      -- CP-element group 623: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Sample/rr
      -- 
    ca_9346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 623_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4156_load_0_ack_1, ack => zeropad3D_CP_2152_elements(623)); -- 
    rr_9359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(623), ack => type_cast_4160_inst_req_0); -- 
    -- CP-element group 624:  transition  input  bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	623 
    -- CP-element group 624: successors 
    -- CP-element group 624:  members (3) 
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_sample_completed_
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Sample/$exit
      -- CP-element group 624: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Sample/ra
      -- 
    ra_9360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4160_inst_ack_0, ack => zeropad3D_CP_2152_elements(624)); -- 
    -- CP-element group 625:  transition  input  bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	620 
    -- CP-element group 625: successors 
    -- CP-element group 625: 	642 
    -- CP-element group 625:  members (3) 
      -- CP-element group 625: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_update_completed_
      -- CP-element group 625: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Update/$exit
      -- CP-element group 625: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4160_Update/ca
      -- 
    ca_9365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4160_inst_ack_1, ack => zeropad3D_CP_2152_elements(625)); -- 
    -- CP-element group 626:  transition  input  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	620 
    -- CP-element group 626: successors 
    -- CP-element group 626:  members (5) 
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_sample_completed_
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/$exit
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/word_access_start/$exit
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/word_access_start/word_0/$exit
      -- CP-element group 626: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Sample/word_access_start/word_0/ra
      -- 
    ra_9382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 626_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4175_load_0_ack_0, ack => zeropad3D_CP_2152_elements(626)); -- 
    -- CP-element group 627:  transition  input  output  bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	620 
    -- CP-element group 627: successors 
    -- CP-element group 627: 	640 
    -- CP-element group 627:  members (12) 
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_update_completed_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/word_access_complete/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/word_access_complete/word_0/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/word_access_complete/word_0/ca
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/LOAD_pad_4175_Merge/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/LOAD_pad_4175_Merge/$exit
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/LOAD_pad_4175_Merge/merge_req
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_pad_4175_Update/LOAD_pad_4175_Merge/merge_ack
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_sample_start_
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Sample/$entry
      -- CP-element group 627: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Sample/rr
      -- 
    ca_9393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4175_load_0_ack_1, ack => zeropad3D_CP_2152_elements(627)); -- 
    rr_9600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(627), ack => type_cast_4252_inst_req_0); -- 
    -- CP-element group 628:  transition  input  bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	620 
    -- CP-element group 628: successors 
    -- CP-element group 628:  members (5) 
      -- CP-element group 628: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_sample_completed_
      -- CP-element group 628: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/$exit
      -- CP-element group 628: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/word_access_start/$exit
      -- CP-element group 628: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/word_access_start/word_0/$exit
      -- CP-element group 628: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Sample/word_access_start/word_0/ra
      -- 
    ra_9415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4178_load_0_ack_0, ack => zeropad3D_CP_2152_elements(628)); -- 
    -- CP-element group 629:  transition  input  output  bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	620 
    -- CP-element group 629: successors 
    -- CP-element group 629: 	636 
    -- CP-element group 629:  members (12) 
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_update_completed_
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/$exit
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/word_access_complete/$exit
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/word_access_complete/word_0/$exit
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/word_access_complete/word_0/ca
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/LOAD_depth_high_4178_Merge/$entry
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/LOAD_depth_high_4178_Merge/$exit
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/LOAD_depth_high_4178_Merge/merge_req
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_depth_high_4178_Update/LOAD_depth_high_4178_Merge/merge_ack
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_sample_start_
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Sample/$entry
      -- CP-element group 629: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Sample/rr
      -- 
    ca_9426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4178_load_0_ack_1, ack => zeropad3D_CP_2152_elements(629)); -- 
    rr_9572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(629), ack => type_cast_4209_inst_req_0); -- 
    -- CP-element group 630:  transition  input  bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	620 
    -- CP-element group 630: successors 
    -- CP-element group 630:  members (5) 
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_sample_completed_
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/$exit
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/word_access_start/$exit
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/word_access_start/word_0/$exit
      -- CP-element group 630: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Sample/word_access_start/word_0/ra
      -- 
    ra_9448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 630_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4181_load_0_ack_0, ack => zeropad3D_CP_2152_elements(630)); -- 
    -- CP-element group 631:  transition  input  output  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	620 
    -- CP-element group 631: successors 
    -- CP-element group 631: 	638 
    -- CP-element group 631:  members (12) 
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_update_completed_
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/$exit
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/word_access_complete/$exit
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/word_access_complete/word_0/$exit
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/word_access_complete/word_0/ca
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/LOAD_col_high_4181_Merge/$entry
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/LOAD_col_high_4181_Merge/$exit
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/LOAD_col_high_4181_Merge/merge_req
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/LOAD_col_high_4181_Update/LOAD_col_high_4181_Merge/merge_ack
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_sample_start_
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Sample/$entry
      -- CP-element group 631: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Sample/rr
      -- 
    ca_9459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 631_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4181_load_0_ack_1, ack => zeropad3D_CP_2152_elements(631)); -- 
    rr_9586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(631), ack => type_cast_4213_inst_req_0); -- 
    -- CP-element group 632:  transition  input  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	620 
    -- CP-element group 632: successors 
    -- CP-element group 632:  members (5) 
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_sample_completed_
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/$exit
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/word_access_start/$exit
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/word_access_start/word_0/$exit
      -- CP-element group 632: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Sample/word_access_start/word_0/ra
      -- 
    ra_9498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4193_load_0_ack_0, ack => zeropad3D_CP_2152_elements(632)); -- 
    -- CP-element group 633:  transition  input  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	620 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	642 
    -- CP-element group 633:  members (9) 
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_update_completed_
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/$exit
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/word_access_complete/$exit
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/word_access_complete/word_0/$exit
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/word_access_complete/word_0/ca
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/ptr_deref_4193_Merge/$entry
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/ptr_deref_4193_Merge/$exit
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/ptr_deref_4193_Merge/merge_req
      -- CP-element group 633: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4193_Update/ptr_deref_4193_Merge/merge_ack
      -- 
    ca_9509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 633_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4193_load_0_ack_1, ack => zeropad3D_CP_2152_elements(633)); -- 
    -- CP-element group 634:  transition  input  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	620 
    -- CP-element group 634: successors 
    -- CP-element group 634:  members (5) 
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_sample_completed_
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/$exit
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/word_access_start/$exit
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/word_access_start/word_0/$exit
      -- CP-element group 634: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Sample/word_access_start/word_0/ra
      -- 
    ra_9548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 634_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4205_load_0_ack_0, ack => zeropad3D_CP_2152_elements(634)); -- 
    -- CP-element group 635:  transition  input  bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	620 
    -- CP-element group 635: successors 
    -- CP-element group 635: 	642 
    -- CP-element group 635:  members (9) 
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_update_completed_
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/word_access_complete/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/word_access_complete/word_0/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/word_access_complete/word_0/ca
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/ptr_deref_4205_Merge/$entry
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/ptr_deref_4205_Merge/$exit
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/ptr_deref_4205_Merge/merge_req
      -- CP-element group 635: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/ptr_deref_4205_Update/ptr_deref_4205_Merge/merge_ack
      -- 
    ca_9559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4205_load_0_ack_1, ack => zeropad3D_CP_2152_elements(635)); -- 
    -- CP-element group 636:  transition  input  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	629 
    -- CP-element group 636: successors 
    -- CP-element group 636:  members (3) 
      -- CP-element group 636: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_sample_completed_
      -- CP-element group 636: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Sample/$exit
      -- CP-element group 636: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Sample/ra
      -- 
    ra_9573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 636_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4209_inst_ack_0, ack => zeropad3D_CP_2152_elements(636)); -- 
    -- CP-element group 637:  transition  input  bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	620 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	642 
    -- CP-element group 637:  members (3) 
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_update_completed_
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Update/$exit
      -- CP-element group 637: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4209_Update/ca
      -- 
    ca_9578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 637_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4209_inst_ack_1, ack => zeropad3D_CP_2152_elements(637)); -- 
    -- CP-element group 638:  transition  input  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	631 
    -- CP-element group 638: successors 
    -- CP-element group 638:  members (3) 
      -- CP-element group 638: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_sample_completed_
      -- CP-element group 638: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Sample/$exit
      -- CP-element group 638: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Sample/ra
      -- 
    ra_9587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 638_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4213_inst_ack_0, ack => zeropad3D_CP_2152_elements(638)); -- 
    -- CP-element group 639:  transition  input  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	620 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	642 
    -- CP-element group 639:  members (3) 
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_update_completed_
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Update/$exit
      -- CP-element group 639: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4213_Update/ca
      -- 
    ca_9592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 639_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4213_inst_ack_1, ack => zeropad3D_CP_2152_elements(639)); -- 
    -- CP-element group 640:  transition  input  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	627 
    -- CP-element group 640: successors 
    -- CP-element group 640:  members (3) 
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_sample_completed_
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Sample/$exit
      -- CP-element group 640: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Sample/ra
      -- 
    ra_9601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4252_inst_ack_0, ack => zeropad3D_CP_2152_elements(640)); -- 
    -- CP-element group 641:  transition  input  bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	620 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	642 
    -- CP-element group 641:  members (3) 
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_update_completed_
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Update/$exit
      -- CP-element group 641: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/type_cast_4252_Update/ca
      -- 
    ca_9606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 641_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4252_inst_ack_1, ack => zeropad3D_CP_2152_elements(641)); -- 
    -- CP-element group 642:  join  fork  transition  place  output  bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	625 
    -- CP-element group 642: 	633 
    -- CP-element group 642: 	635 
    -- CP-element group 642: 	637 
    -- CP-element group 642: 	639 
    -- CP-element group 642: 	641 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	1108 
    -- CP-element group 642: 	1109 
    -- CP-element group 642: 	1110 
    -- CP-element group 642: 	1112 
    -- CP-element group 642:  members (16) 
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341
      -- CP-element group 642: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294__exit__
      -- CP-element group 642: 	 branch_block_stmt_714/assign_stmt_4157_to_assign_stmt_4294/$exit
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4310/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Update/cr
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Update/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Sample/rr
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Sample/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4297/$entry
      -- CP-element group 642: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/$entry
      -- 
    cr_13807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(642), ack => type_cast_4307_inst_req_1); -- 
    rr_13802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(642), ack => type_cast_4307_inst_req_0); -- 
    zeropad3D_cp_element_group_642: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_642"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(625) & zeropad3D_CP_2152_elements(633) & zeropad3D_CP_2152_elements(635) & zeropad3D_CP_2152_elements(637) & zeropad3D_CP_2152_elements(639) & zeropad3D_CP_2152_elements(641);
      gj_zeropad3D_cp_element_group_642 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(642), clk => clk, reset => reset); --
    end block;
    -- CP-element group 643:  transition  input  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	1118 
    -- CP-element group 643: successors 
    -- CP-element group 643:  members (3) 
      -- CP-element group 643: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_sample_completed_
      -- CP-element group 643: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Sample/$exit
      -- CP-element group 643: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Sample/ra
      -- 
    ra_9618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 643_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4321_inst_ack_0, ack => zeropad3D_CP_2152_elements(643)); -- 
    -- CP-element group 644:  branch  transition  place  input  output  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	1118 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644: 	646 
    -- CP-element group 644:  members (13) 
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330__entry__
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329__exit__
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/$exit
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_update_completed_
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Update/$exit
      -- CP-element group 644: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Update/ca
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330_dead_link/$entry
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330_eval_test/$entry
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330_eval_test/$exit
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330_eval_test/branch_req
      -- CP-element group 644: 	 branch_block_stmt_714/R_cmp1346_4331_place
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330_if_link/$entry
      -- CP-element group 644: 	 branch_block_stmt_714/if_stmt_4330_else_link/$entry
      -- 
    ca_9623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 644_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4321_inst_ack_1, ack => zeropad3D_CP_2152_elements(644)); -- 
    branch_req_9631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(644), ack => if_stmt_4330_branch_req_0); -- 
    -- CP-element group 645:  transition  place  input  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645: 	1119 
    -- CP-element group 645:  members (5) 
      -- CP-element group 645: 	 branch_block_stmt_714/if_stmt_4330_if_link/$exit
      -- CP-element group 645: 	 branch_block_stmt_714/if_stmt_4330_if_link/if_choice_transition
      -- CP-element group 645: 	 branch_block_stmt_714/whilex_xbody1341_ifx_xthen1376
      -- CP-element group 645: 	 branch_block_stmt_714/whilex_xbody1341_ifx_xthen1376_PhiReq/$exit
      -- CP-element group 645: 	 branch_block_stmt_714/whilex_xbody1341_ifx_xthen1376_PhiReq/$entry
      -- 
    if_choice_transition_9636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 645_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4330_branch_ack_1, ack => zeropad3D_CP_2152_elements(645)); -- 
    -- CP-element group 646:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	644 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	647 
    -- CP-element group 646: 	648 
    -- CP-element group 646: 	650 
    -- CP-element group 646:  members (27) 
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355__entry__
      -- CP-element group 646: 	 branch_block_stmt_714/merge_stmt_4336__exit__
      -- CP-element group 646: 	 branch_block_stmt_714/if_stmt_4330_else_link/$exit
      -- CP-element group 646: 	 branch_block_stmt_714/if_stmt_4330_else_link/else_choice_transition
      -- CP-element group 646: 	 branch_block_stmt_714/whilex_xbody1341_lorx_xlhsx_xfalse1348
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_sample_start_
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_update_start_
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_word_address_calculated
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_root_address_calculated
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/word_access_start/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/word_access_start/word_0/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/word_access_start/word_0/rr
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/word_access_complete/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/word_access_complete/word_0/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/word_access_complete/word_0/cr
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_update_start_
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Update/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Update/cr
      -- CP-element group 646: 	 branch_block_stmt_714/whilex_xbody1341_lorx_xlhsx_xfalse1348_PhiReq/$exit
      -- CP-element group 646: 	 branch_block_stmt_714/merge_stmt_4336_PhiAck/$entry
      -- CP-element group 646: 	 branch_block_stmt_714/merge_stmt_4336_PhiAck/$exit
      -- CP-element group 646: 	 branch_block_stmt_714/merge_stmt_4336_PhiAck/dummy
      -- CP-element group 646: 	 branch_block_stmt_714/merge_stmt_4336_PhiReqMerge
      -- CP-element group 646: 	 branch_block_stmt_714/whilex_xbody1341_lorx_xlhsx_xfalse1348_PhiReq/$entry
      -- 
    else_choice_transition_9640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 646_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4330_branch_ack_0, ack => zeropad3D_CP_2152_elements(646)); -- 
    rr_9661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(646), ack => LOAD_row_high_4338_load_0_req_0); -- 
    cr_9672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(646), ack => LOAD_row_high_4338_load_0_req_1); -- 
    cr_9691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(646), ack => type_cast_4342_inst_req_1); -- 
    -- CP-element group 647:  transition  input  bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	646 
    -- CP-element group 647: successors 
    -- CP-element group 647:  members (5) 
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_sample_completed_
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/$exit
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/word_access_start/$exit
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/word_access_start/word_0/$exit
      -- CP-element group 647: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Sample/word_access_start/word_0/ra
      -- 
    ra_9662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4338_load_0_ack_0, ack => zeropad3D_CP_2152_elements(647)); -- 
    -- CP-element group 648:  transition  input  output  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	646 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (12) 
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_update_completed_
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/$exit
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/word_access_complete/$exit
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/word_access_complete/word_0/$exit
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/word_access_complete/word_0/ca
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/LOAD_row_high_4338_Merge/$entry
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/LOAD_row_high_4338_Merge/$exit
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/LOAD_row_high_4338_Merge/merge_req
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/LOAD_row_high_4338_Update/LOAD_row_high_4338_Merge/merge_ack
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_sample_start_
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Sample/$entry
      -- CP-element group 648: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Sample/rr
      -- 
    ca_9673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 648_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4338_load_0_ack_1, ack => zeropad3D_CP_2152_elements(648)); -- 
    rr_9686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(648), ack => type_cast_4342_inst_req_0); -- 
    -- CP-element group 649:  transition  input  bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649:  members (3) 
      -- CP-element group 649: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_sample_completed_
      -- CP-element group 649: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Sample/$exit
      -- CP-element group 649: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Sample/ra
      -- 
    ra_9687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 649_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4342_inst_ack_0, ack => zeropad3D_CP_2152_elements(649)); -- 
    -- CP-element group 650:  branch  transition  place  input  output  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	646 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	651 
    -- CP-element group 650: 	652 
    -- CP-element group 650:  members (13) 
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355__exit__
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356__entry__
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_update_completed_
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Update/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/assign_stmt_4339_to_assign_stmt_4355/type_cast_4342_Update/ca
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356_dead_link/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356_eval_test/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356_eval_test/$exit
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356_eval_test/branch_req
      -- CP-element group 650: 	 branch_block_stmt_714/R_cmp1356_4357_place
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356_if_link/$entry
      -- CP-element group 650: 	 branch_block_stmt_714/if_stmt_4356_else_link/$entry
      -- 
    ca_9692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 650_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4342_inst_ack_1, ack => zeropad3D_CP_2152_elements(650)); -- 
    branch_req_9700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(650), ack => if_stmt_4356_branch_req_0); -- 
    -- CP-element group 651:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	650 
    -- CP-element group 651: successors 
    -- CP-element group 651: 	653 
    -- CP-element group 651: 	654 
    -- CP-element group 651:  members (18) 
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374__entry__
      -- CP-element group 651: 	 branch_block_stmt_714/merge_stmt_4362__exit__
      -- CP-element group 651: 	 branch_block_stmt_714/if_stmt_4356_if_link/$exit
      -- CP-element group 651: 	 branch_block_stmt_714/if_stmt_4356_if_link/if_choice_transition
      -- CP-element group 651: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1358
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/$entry
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_sample_start_
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_update_start_
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Sample/$entry
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Sample/rr
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Update/$entry
      -- CP-element group 651: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Update/cr
      -- CP-element group 651: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1358_PhiReq/$entry
      -- CP-element group 651: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_lorx_xlhsx_xfalse1358_PhiReq/$exit
      -- CP-element group 651: 	 branch_block_stmt_714/merge_stmt_4362_PhiReqMerge
      -- CP-element group 651: 	 branch_block_stmt_714/merge_stmt_4362_PhiAck/$entry
      -- CP-element group 651: 	 branch_block_stmt_714/merge_stmt_4362_PhiAck/$exit
      -- CP-element group 651: 	 branch_block_stmt_714/merge_stmt_4362_PhiAck/dummy
      -- 
    if_choice_transition_9705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 651_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4356_branch_ack_1, ack => zeropad3D_CP_2152_elements(651)); -- 
    rr_9722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(651), ack => type_cast_4366_inst_req_0); -- 
    cr_9727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(651), ack => type_cast_4366_inst_req_1); -- 
    -- CP-element group 652:  transition  place  input  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	650 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	1119 
    -- CP-element group 652:  members (5) 
      -- CP-element group 652: 	 branch_block_stmt_714/if_stmt_4356_else_link/$exit
      -- CP-element group 652: 	 branch_block_stmt_714/if_stmt_4356_else_link/else_choice_transition
      -- CP-element group 652: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_ifx_xthen1376
      -- CP-element group 652: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_ifx_xthen1376_PhiReq/$exit
      -- CP-element group 652: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1348_ifx_xthen1376_PhiReq/$entry
      -- 
    else_choice_transition_9709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4356_branch_ack_0, ack => zeropad3D_CP_2152_elements(652)); -- 
    -- CP-element group 653:  transition  input  bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	651 
    -- CP-element group 653: successors 
    -- CP-element group 653:  members (3) 
      -- CP-element group 653: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_sample_completed_
      -- CP-element group 653: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Sample/$exit
      -- CP-element group 653: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Sample/ra
      -- 
    ra_9723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 653_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4366_inst_ack_0, ack => zeropad3D_CP_2152_elements(653)); -- 
    -- CP-element group 654:  branch  transition  place  input  output  bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	651 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	655 
    -- CP-element group 654: 	656 
    -- CP-element group 654:  members (13) 
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374__exit__
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375__entry__
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/$exit
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_update_completed_
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Update/$exit
      -- CP-element group 654: 	 branch_block_stmt_714/assign_stmt_4367_to_assign_stmt_4374/type_cast_4366_Update/ca
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375_dead_link/$entry
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375_eval_test/$entry
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375_eval_test/$exit
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375_eval_test/branch_req
      -- CP-element group 654: 	 branch_block_stmt_714/R_cmp1363_4376_place
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375_if_link/$entry
      -- CP-element group 654: 	 branch_block_stmt_714/if_stmt_4375_else_link/$entry
      -- 
    ca_9728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 654_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4366_inst_ack_1, ack => zeropad3D_CP_2152_elements(654)); -- 
    branch_req_9736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(654), ack => if_stmt_4375_branch_req_0); -- 
    -- CP-element group 655:  transition  place  input  bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	654 
    -- CP-element group 655: successors 
    -- CP-element group 655: 	1119 
    -- CP-element group 655:  members (5) 
      -- CP-element group 655: 	 branch_block_stmt_714/if_stmt_4375_if_link/$exit
      -- CP-element group 655: 	 branch_block_stmt_714/if_stmt_4375_if_link/if_choice_transition
      -- CP-element group 655: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_ifx_xthen1376
      -- CP-element group 655: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_ifx_xthen1376_PhiReq/$exit
      -- CP-element group 655: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_ifx_xthen1376_PhiReq/$entry
      -- 
    if_choice_transition_9741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4375_branch_ack_1, ack => zeropad3D_CP_2152_elements(655)); -- 
    -- CP-element group 656:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	654 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	657 
    -- CP-element group 656: 	658 
    -- CP-element group 656: 	660 
    -- CP-element group 656:  members (27) 
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406__entry__
      -- CP-element group 656: 	 branch_block_stmt_714/merge_stmt_4381__exit__
      -- CP-element group 656: 	 branch_block_stmt_714/if_stmt_4375_else_link/$exit
      -- CP-element group 656: 	 branch_block_stmt_714/if_stmt_4375_else_link/else_choice_transition
      -- CP-element group 656: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_lorx_xlhsx_xfalse1365
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_sample_start_
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_update_start_
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_word_address_calculated
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_root_address_calculated
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/word_access_start/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/word_access_start/word_0/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/word_access_start/word_0/rr
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/word_access_complete/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/word_access_complete/word_0/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/word_access_complete/word_0/cr
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_update_start_
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Update/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Update/cr
      -- CP-element group 656: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_lorx_xlhsx_xfalse1365_PhiReq/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1358_lorx_xlhsx_xfalse1365_PhiReq/$exit
      -- CP-element group 656: 	 branch_block_stmt_714/merge_stmt_4381_PhiReqMerge
      -- CP-element group 656: 	 branch_block_stmt_714/merge_stmt_4381_PhiAck/$entry
      -- CP-element group 656: 	 branch_block_stmt_714/merge_stmt_4381_PhiAck/$exit
      -- CP-element group 656: 	 branch_block_stmt_714/merge_stmt_4381_PhiAck/dummy
      -- 
    else_choice_transition_9745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4375_branch_ack_0, ack => zeropad3D_CP_2152_elements(656)); -- 
    rr_9766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(656), ack => LOAD_col_high_4383_load_0_req_0); -- 
    cr_9777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(656), ack => LOAD_col_high_4383_load_0_req_1); -- 
    cr_9796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(656), ack => type_cast_4387_inst_req_1); -- 
    -- CP-element group 657:  transition  input  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	656 
    -- CP-element group 657: successors 
    -- CP-element group 657:  members (5) 
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_sample_completed_
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/$exit
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/word_access_start/$exit
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/word_access_start/word_0/$exit
      -- CP-element group 657: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Sample/word_access_start/word_0/ra
      -- 
    ra_9767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 657_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4383_load_0_ack_0, ack => zeropad3D_CP_2152_elements(657)); -- 
    -- CP-element group 658:  transition  input  output  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	656 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	659 
    -- CP-element group 658:  members (12) 
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_update_completed_
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/word_access_complete/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/word_access_complete/word_0/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/word_access_complete/word_0/ca
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/LOAD_col_high_4383_Merge/$entry
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/LOAD_col_high_4383_Merge/$exit
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/LOAD_col_high_4383_Merge/merge_req
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/LOAD_col_high_4383_Update/LOAD_col_high_4383_Merge/merge_ack
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_sample_start_
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Sample/$entry
      -- CP-element group 658: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Sample/rr
      -- 
    ca_9778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 658_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4383_load_0_ack_1, ack => zeropad3D_CP_2152_elements(658)); -- 
    rr_9791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(658), ack => type_cast_4387_inst_req_0); -- 
    -- CP-element group 659:  transition  input  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	658 
    -- CP-element group 659: successors 
    -- CP-element group 659:  members (3) 
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_sample_completed_
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Sample/$exit
      -- CP-element group 659: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Sample/ra
      -- 
    ra_9792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 659_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4387_inst_ack_0, ack => zeropad3D_CP_2152_elements(659)); -- 
    -- CP-element group 660:  branch  transition  place  input  output  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	656 
    -- CP-element group 660: successors 
    -- CP-element group 660: 	661 
    -- CP-element group 660: 	662 
    -- CP-element group 660:  members (13) 
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406__exit__
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407__entry__
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/$exit
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_update_completed_
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Update/$exit
      -- CP-element group 660: 	 branch_block_stmt_714/assign_stmt_4384_to_assign_stmt_4406/type_cast_4387_Update/ca
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407_dead_link/$entry
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407_eval_test/$entry
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407_eval_test/$exit
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407_eval_test/branch_req
      -- CP-element group 660: 	 branch_block_stmt_714/R_cmp1374_4408_place
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407_if_link/$entry
      -- CP-element group 660: 	 branch_block_stmt_714/if_stmt_4407_else_link/$entry
      -- 
    ca_9797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4387_inst_ack_1, ack => zeropad3D_CP_2152_elements(660)); -- 
    branch_req_9805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(660), ack => if_stmt_4407_branch_req_0); -- 
    -- CP-element group 661:  fork  transition  place  input  output  bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	660 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	677 
    -- CP-element group 661: 	678 
    -- CP-element group 661: 	680 
    -- CP-element group 661: 	682 
    -- CP-element group 661: 	684 
    -- CP-element group 661: 	686 
    -- CP-element group 661: 	688 
    -- CP-element group 661: 	690 
    -- CP-element group 661: 	692 
    -- CP-element group 661: 	695 
    -- CP-element group 661:  members (46) 
      -- CP-element group 661: 	 branch_block_stmt_714/merge_stmt_4471__exit__
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576__entry__
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/word_access_complete/word_0/cr
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_complete/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_complete/req
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Update/cr
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Update/req
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/word_access_complete/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/word_access_complete/word_0/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_update_start
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/word_access_complete/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/word_access_complete/word_0/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/word_access_complete/word_0/cr
      -- CP-element group 661: 	 branch_block_stmt_714/if_stmt_4407_if_link/$exit
      -- CP-element group 661: 	 branch_block_stmt_714/if_stmt_4407_if_link/if_choice_transition
      -- CP-element group 661: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xelse1397
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_sample_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Sample/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Sample/rr
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Update/cr
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Update/cr
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_update_start
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Update/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Update/req
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_complete/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_complete/req
      -- CP-element group 661: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_update_start_
      -- CP-element group 661: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xelse1397_PhiReq/$entry
      -- CP-element group 661: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xelse1397_PhiReq/$exit
      -- CP-element group 661: 	 branch_block_stmt_714/merge_stmt_4471_PhiReqMerge
      -- CP-element group 661: 	 branch_block_stmt_714/merge_stmt_4471_PhiAck/dummy
      -- CP-element group 661: 	 branch_block_stmt_714/merge_stmt_4471_PhiAck/$exit
      -- CP-element group 661: 	 branch_block_stmt_714/merge_stmt_4471_PhiAck/$entry
      -- 
    if_choice_transition_9810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 661_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4407_branch_ack_1, ack => zeropad3D_CP_2152_elements(661)); -- 
    cr_10193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => ptr_deref_4574_store_0_req_1); -- 
    req_10143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => addr_of_4571_final_reg_req_1); -- 
    cr_10097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => type_cast_4564_inst_req_1); -- 
    req_10128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => array_obj_ref_4570_index_offset_req_1); -- 
    cr_10078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => ptr_deref_4550_load_0_req_1); -- 
    rr_9968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => type_cast_4475_inst_req_0); -- 
    cr_9973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => type_cast_4475_inst_req_1); -- 
    cr_9987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => type_cast_4539_inst_req_1); -- 
    req_10018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => array_obj_ref_4545_index_offset_req_1); -- 
    req_10033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(661), ack => addr_of_4546_final_reg_req_1); -- 
    -- CP-element group 662:  transition  place  input  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	660 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	1119 
    -- CP-element group 662:  members (5) 
      -- CP-element group 662: 	 branch_block_stmt_714/if_stmt_4407_else_link/$exit
      -- CP-element group 662: 	 branch_block_stmt_714/if_stmt_4407_else_link/else_choice_transition
      -- CP-element group 662: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xthen1376
      -- CP-element group 662: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xthen1376_PhiReq/$exit
      -- CP-element group 662: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1365_ifx_xthen1376_PhiReq/$entry
      -- 
    else_choice_transition_9814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 662_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4407_branch_ack_0, ack => zeropad3D_CP_2152_elements(662)); -- 
    -- CP-element group 663:  transition  input  bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	1119 
    -- CP-element group 663: successors 
    -- CP-element group 663:  members (3) 
      -- CP-element group 663: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_sample_completed_
      -- CP-element group 663: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Sample/$exit
      -- CP-element group 663: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Sample/ra
      -- 
    ra_9828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4417_inst_ack_0, ack => zeropad3D_CP_2152_elements(663)); -- 
    -- CP-element group 664:  transition  input  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	1119 
    -- CP-element group 664: successors 
    -- CP-element group 664: 	667 
    -- CP-element group 664:  members (3) 
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_update_completed_
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Update/$exit
      -- CP-element group 664: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Update/ca
      -- 
    ca_9833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 664_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4417_inst_ack_1, ack => zeropad3D_CP_2152_elements(664)); -- 
    -- CP-element group 665:  transition  input  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	1119 
    -- CP-element group 665: successors 
    -- CP-element group 665:  members (3) 
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_sample_completed_
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Sample/$exit
      -- CP-element group 665: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Sample/ra
      -- 
    ra_9842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 665_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4422_inst_ack_0, ack => zeropad3D_CP_2152_elements(665)); -- 
    -- CP-element group 666:  transition  input  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	1119 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	667 
    -- CP-element group 666:  members (3) 
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_update_completed_
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Update/$exit
      -- CP-element group 666: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Update/ca
      -- 
    ca_9847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 666_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4422_inst_ack_1, ack => zeropad3D_CP_2152_elements(666)); -- 
    -- CP-element group 667:  join  transition  output  bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	664 
    -- CP-element group 667: 	666 
    -- CP-element group 667: successors 
    -- CP-element group 667: 	668 
    -- CP-element group 667:  members (3) 
      -- CP-element group 667: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_sample_start_
      -- CP-element group 667: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Sample/$entry
      -- CP-element group 667: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Sample/rr
      -- 
    rr_9855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(667), ack => type_cast_4456_inst_req_0); -- 
    zeropad3D_cp_element_group_667: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_667"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(664) & zeropad3D_CP_2152_elements(666);
      gj_zeropad3D_cp_element_group_667 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(667), clk => clk, reset => reset); --
    end block;
    -- CP-element group 668:  transition  input  bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	667 
    -- CP-element group 668: successors 
    -- CP-element group 668:  members (3) 
      -- CP-element group 668: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_sample_completed_
      -- CP-element group 668: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Sample/$exit
      -- CP-element group 668: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Sample/ra
      -- 
    ra_9856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 668_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4456_inst_ack_0, ack => zeropad3D_CP_2152_elements(668)); -- 
    -- CP-element group 669:  transition  input  output  bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	1119 
    -- CP-element group 669: successors 
    -- CP-element group 669: 	670 
    -- CP-element group 669:  members (16) 
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_update_completed_
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Update/$exit
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Update/ca
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_resized_1
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_scaled_1
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_computed_1
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_resize_1/$entry
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_resize_1/$exit
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_resize_1/index_resize_req
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_resize_1/index_resize_ack
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_scale_1/$entry
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_scale_1/$exit
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_scale_1/scale_rename_req
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_index_scale_1/scale_rename_ack
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Sample/$entry
      -- CP-element group 669: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Sample/req
      -- 
    ca_9861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 669_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4456_inst_ack_1, ack => zeropad3D_CP_2152_elements(669)); -- 
    req_9886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(669), ack => array_obj_ref_4462_index_offset_req_0); -- 
    -- CP-element group 670:  transition  input  bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	669 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	676 
    -- CP-element group 670:  members (3) 
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_sample_complete
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Sample/$exit
      -- CP-element group 670: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Sample/ack
      -- 
    ack_9887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 670_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4462_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(670)); -- 
    -- CP-element group 671:  transition  input  output  bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	1119 
    -- CP-element group 671: successors 
    -- CP-element group 671: 	672 
    -- CP-element group 671:  members (11) 
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_sample_start_
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_root_address_calculated
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_offset_calculated
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Update/$exit
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Update/ack
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_base_plus_offset/$entry
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_base_plus_offset/$exit
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_base_plus_offset/sum_rename_req
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_base_plus_offset/sum_rename_ack
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_request/$entry
      -- CP-element group 671: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_request/req
      -- 
    ack_9892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4462_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(671)); -- 
    req_9901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(671), ack => addr_of_4463_final_reg_req_0); -- 
    -- CP-element group 672:  transition  input  bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	671 
    -- CP-element group 672: successors 
    -- CP-element group 672:  members (3) 
      -- CP-element group 672: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_sample_completed_
      -- CP-element group 672: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_request/$exit
      -- CP-element group 672: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_request/ack
      -- 
    ack_9902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4463_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(672)); -- 
    -- CP-element group 673:  join  fork  transition  input  output  bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	1119 
    -- CP-element group 673: successors 
    -- CP-element group 673: 	674 
    -- CP-element group 673:  members (28) 
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_update_completed_
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_complete/$exit
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_complete/ack
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_sample_start_
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_address_calculated
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_word_address_calculated
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_root_address_calculated
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_address_resized
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_addr_resize/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_addr_resize/$exit
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_addr_resize/base_resize_req
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_addr_resize/base_resize_ack
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_plus_offset/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_plus_offset/$exit
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_plus_offset/sum_rename_req
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_base_plus_offset/sum_rename_ack
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_word_addrgen/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_word_addrgen/$exit
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_word_addrgen/root_register_req
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_word_addrgen/root_register_ack
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/ptr_deref_4466_Split/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/ptr_deref_4466_Split/$exit
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/ptr_deref_4466_Split/split_req
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/ptr_deref_4466_Split/split_ack
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/word_access_start/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/word_access_start/word_0/$entry
      -- CP-element group 673: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/word_access_start/word_0/rr
      -- 
    ack_9907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 673_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4463_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(673)); -- 
    rr_9945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(673), ack => ptr_deref_4466_store_0_req_0); -- 
    -- CP-element group 674:  transition  input  bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	673 
    -- CP-element group 674: successors 
    -- CP-element group 674:  members (5) 
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_sample_completed_
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/$exit
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/word_access_start/$exit
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/word_access_start/word_0/$exit
      -- CP-element group 674: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Sample/word_access_start/word_0/ra
      -- 
    ra_9946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 674_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4466_store_0_ack_0, ack => zeropad3D_CP_2152_elements(674)); -- 
    -- CP-element group 675:  transition  input  bypass 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	1119 
    -- CP-element group 675: successors 
    -- CP-element group 675: 	676 
    -- CP-element group 675:  members (5) 
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_update_completed_
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/$exit
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/word_access_complete/$exit
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/word_access_complete/word_0/$exit
      -- CP-element group 675: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/word_access_complete/word_0/ca
      -- 
    ca_9957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4466_store_0_ack_1, ack => zeropad3D_CP_2152_elements(675)); -- 
    -- CP-element group 676:  join  transition  place  bypass 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	670 
    -- CP-element group 676: 	675 
    -- CP-element group 676: successors 
    -- CP-element group 676: 	1120 
    -- CP-element group 676:  members (5) 
      -- CP-element group 676: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469__exit__
      -- CP-element group 676: 	 branch_block_stmt_714/ifx_xthen1376_ifx_xend1445
      -- CP-element group 676: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/$exit
      -- CP-element group 676: 	 branch_block_stmt_714/ifx_xthen1376_ifx_xend1445_PhiReq/$exit
      -- CP-element group 676: 	 branch_block_stmt_714/ifx_xthen1376_ifx_xend1445_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_676: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_676"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(670) & zeropad3D_CP_2152_elements(675);
      gj_zeropad3D_cp_element_group_676 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(676), clk => clk, reset => reset); --
    end block;
    -- CP-element group 677:  transition  input  bypass 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	661 
    -- CP-element group 677: successors 
    -- CP-element group 677:  members (3) 
      -- CP-element group 677: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_sample_completed_
      -- CP-element group 677: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Sample/$exit
      -- CP-element group 677: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Sample/ra
      -- 
    ra_9969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 677_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4475_inst_ack_0, ack => zeropad3D_CP_2152_elements(677)); -- 
    -- CP-element group 678:  fork  transition  input  output  bypass 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: 	661 
    -- CP-element group 678: successors 
    -- CP-element group 678: 	679 
    -- CP-element group 678: 	687 
    -- CP-element group 678:  members (9) 
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Sample/rr
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Sample/$entry
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_sample_start_
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_update_completed_
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Update/$exit
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4475_Update/ca
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_sample_start_
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Sample/$entry
      -- CP-element group 678: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Sample/rr
      -- 
    ca_9974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 678_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4475_inst_ack_1, ack => zeropad3D_CP_2152_elements(678)); -- 
    rr_9982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(678), ack => type_cast_4539_inst_req_0); -- 
    rr_10092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(678), ack => type_cast_4564_inst_req_0); -- 
    -- CP-element group 679:  transition  input  bypass 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	678 
    -- CP-element group 679: successors 
    -- CP-element group 679:  members (3) 
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_sample_completed_
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Sample/$exit
      -- CP-element group 679: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Sample/ra
      -- 
    ra_9983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 679_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4539_inst_ack_0, ack => zeropad3D_CP_2152_elements(679)); -- 
    -- CP-element group 680:  transition  input  output  bypass 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	661 
    -- CP-element group 680: successors 
    -- CP-element group 680: 	681 
    -- CP-element group 680:  members (16) 
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_update_completed_
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Update/$exit
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4539_Update/ca
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_resized_1
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_scaled_1
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_computed_1
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_resize_1/$entry
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_resize_1/$exit
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_resize_1/index_resize_req
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_resize_1/index_resize_ack
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_scale_1/$entry
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_scale_1/$exit
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_scale_1/scale_rename_req
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_index_scale_1/scale_rename_ack
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Sample/$entry
      -- CP-element group 680: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Sample/req
      -- 
    ca_9988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 680_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4539_inst_ack_1, ack => zeropad3D_CP_2152_elements(680)); -- 
    req_10013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(680), ack => array_obj_ref_4545_index_offset_req_0); -- 
    -- CP-element group 681:  transition  input  bypass 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	680 
    -- CP-element group 681: successors 
    -- CP-element group 681: 	696 
    -- CP-element group 681:  members (3) 
      -- CP-element group 681: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_sample_complete
      -- CP-element group 681: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Sample/$exit
      -- CP-element group 681: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Sample/ack
      -- 
    ack_10014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 681_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4545_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(681)); -- 
    -- CP-element group 682:  transition  input  output  bypass 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	661 
    -- CP-element group 682: successors 
    -- CP-element group 682: 	683 
    -- CP-element group 682:  members (11) 
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_sample_start_
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_root_address_calculated
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_offset_calculated
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Update/$exit
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_final_index_sum_regn_Update/ack
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_base_plus_offset/$entry
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_base_plus_offset/$exit
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_base_plus_offset/sum_rename_req
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4545_base_plus_offset/sum_rename_ack
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_request/$entry
      -- CP-element group 682: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_request/req
      -- 
    ack_10019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 682_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4545_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(682)); -- 
    req_10028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(682), ack => addr_of_4546_final_reg_req_0); -- 
    -- CP-element group 683:  transition  input  bypass 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	682 
    -- CP-element group 683: successors 
    -- CP-element group 683:  members (3) 
      -- CP-element group 683: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_sample_completed_
      -- CP-element group 683: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_request/$exit
      -- CP-element group 683: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_request/ack
      -- 
    ack_10029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 683_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4546_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(683)); -- 
    -- CP-element group 684:  join  fork  transition  input  output  bypass 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	661 
    -- CP-element group 684: successors 
    -- CP-element group 684: 	685 
    -- CP-element group 684:  members (24) 
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/word_access_start/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/word_access_start/word_0/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/word_access_start/word_0/rr
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_update_completed_
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_complete/$exit
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4546_complete/ack
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_sample_start_
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_address_calculated
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_word_address_calculated
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_root_address_calculated
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_address_resized
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_addr_resize/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_addr_resize/$exit
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_addr_resize/base_resize_req
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_addr_resize/base_resize_ack
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_plus_offset/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_plus_offset/$exit
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_plus_offset/sum_rename_req
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_base_plus_offset/sum_rename_ack
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_word_addrgen/$entry
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_word_addrgen/$exit
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_word_addrgen/root_register_req
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_word_addrgen/root_register_ack
      -- CP-element group 684: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/$entry
      -- 
    ack_10034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 684_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4546_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(684)); -- 
    rr_10067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(684), ack => ptr_deref_4550_load_0_req_0); -- 
    -- CP-element group 685:  transition  input  bypass 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	684 
    -- CP-element group 685: successors 
    -- CP-element group 685:  members (5) 
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/word_access_start/$exit
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/word_access_start/word_0/$exit
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/word_access_start/word_0/ra
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_sample_completed_
      -- CP-element group 685: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Sample/$exit
      -- 
    ra_10068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 685_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4550_load_0_ack_0, ack => zeropad3D_CP_2152_elements(685)); -- 
    -- CP-element group 686:  transition  input  bypass 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: 	661 
    -- CP-element group 686: successors 
    -- CP-element group 686: 	693 
    -- CP-element group 686:  members (9) 
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/$exit
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/word_access_complete/$exit
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/ptr_deref_4550_Merge/merge_ack
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/ptr_deref_4550_Merge/merge_req
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/ptr_deref_4550_Merge/$exit
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/ptr_deref_4550_Merge/$entry
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/word_access_complete/word_0/ca
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_Update/word_access_complete/word_0/$exit
      -- CP-element group 686: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4550_update_completed_
      -- 
    ca_10079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 686_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4550_load_0_ack_1, ack => zeropad3D_CP_2152_elements(686)); -- 
    -- CP-element group 687:  transition  input  bypass 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	678 
    -- CP-element group 687: successors 
    -- CP-element group 687:  members (3) 
      -- CP-element group 687: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Sample/$exit
      -- CP-element group 687: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Sample/ra
      -- CP-element group 687: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_sample_completed_
      -- 
    ra_10093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4564_inst_ack_0, ack => zeropad3D_CP_2152_elements(687)); -- 
    -- CP-element group 688:  transition  input  output  bypass 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	661 
    -- CP-element group 688: successors 
    -- CP-element group 688: 	689 
    -- CP-element group 688:  members (16) 
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_computed_1
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_resize_1/$entry
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_resize_1/$exit
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_resize_1/index_resize_req
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_resize_1/index_resize_ack
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Update/$exit
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_Update/ca
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_scale_1/$entry
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_scale_1/$exit
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_scale_1/scale_rename_req
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_scale_1/scale_rename_ack
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Sample/$entry
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Sample/req
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_resized_1
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_index_scaled_1
      -- CP-element group 688: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/type_cast_4564_update_completed_
      -- 
    ca_10098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 688_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4564_inst_ack_1, ack => zeropad3D_CP_2152_elements(688)); -- 
    req_10123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(688), ack => array_obj_ref_4570_index_offset_req_0); -- 
    -- CP-element group 689:  transition  input  bypass 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	688 
    -- CP-element group 689: successors 
    -- CP-element group 689: 	696 
    -- CP-element group 689:  members (3) 
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_sample_complete
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Sample/$exit
      -- CP-element group 689: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Sample/ack
      -- 
    ack_10124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 689_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4570_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(689)); -- 
    -- CP-element group 690:  transition  input  output  bypass 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	661 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	691 
    -- CP-element group 690:  members (11) 
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_base_plus_offset/sum_rename_ack
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_request/$entry
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_request/req
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Update/$exit
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_final_index_sum_regn_Update/ack
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_base_plus_offset/$entry
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_sample_start_
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_root_address_calculated
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_base_plus_offset/$exit
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_offset_calculated
      -- CP-element group 690: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/array_obj_ref_4570_base_plus_offset/sum_rename_req
      -- 
    ack_10129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 690_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_4570_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(690)); -- 
    req_10138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(690), ack => addr_of_4571_final_reg_req_0); -- 
    -- CP-element group 691:  transition  input  bypass 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	690 
    -- CP-element group 691: successors 
    -- CP-element group 691:  members (3) 
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_request/$exit
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_request/ack
      -- CP-element group 691: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_sample_completed_
      -- 
    ack_10139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 691_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4571_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(691)); -- 
    -- CP-element group 692:  fork  transition  input  bypass 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	661 
    -- CP-element group 692: successors 
    -- CP-element group 692: 	693 
    -- CP-element group 692:  members (19) 
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_addr_resize/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_complete/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_addr_resize/base_resize_req
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_complete/ack
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/addr_of_4571_update_completed_
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_addr_resize/base_resize_ack
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_plus_offset/$entry
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_address_calculated
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_word_address_calculated
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_root_address_calculated
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_address_resized
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_plus_offset/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_plus_offset/sum_rename_req
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_addr_resize/$entry
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_base_plus_offset/sum_rename_ack
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_word_addrgen/root_register_ack
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_word_addrgen/root_register_req
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_word_addrgen/$exit
      -- CP-element group 692: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_word_addrgen/$entry
      -- 
    ack_10144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_4571_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(692)); -- 
    -- CP-element group 693:  join  transition  output  bypass 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	686 
    -- CP-element group 693: 	692 
    -- CP-element group 693: successors 
    -- CP-element group 693: 	694 
    -- CP-element group 693:  members (9) 
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/$entry
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/ptr_deref_4574_Split/$entry
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/ptr_deref_4574_Split/$exit
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/ptr_deref_4574_Split/split_req
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/ptr_deref_4574_Split/split_ack
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/word_access_start/$entry
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_sample_start_
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/word_access_start/word_0/$entry
      -- CP-element group 693: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/word_access_start/word_0/rr
      -- 
    rr_10182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(693), ack => ptr_deref_4574_store_0_req_0); -- 
    zeropad3D_cp_element_group_693: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_693"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(686) & zeropad3D_CP_2152_elements(692);
      gj_zeropad3D_cp_element_group_693 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(693), clk => clk, reset => reset); --
    end block;
    -- CP-element group 694:  transition  input  bypass 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	693 
    -- CP-element group 694: successors 
    -- CP-element group 694:  members (5) 
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/$exit
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/word_access_start/$exit
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/word_access_start/word_0/$exit
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_sample_completed_
      -- CP-element group 694: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Sample/word_access_start/word_0/ra
      -- 
    ra_10183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 694_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4574_store_0_ack_0, ack => zeropad3D_CP_2152_elements(694)); -- 
    -- CP-element group 695:  transition  input  bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	661 
    -- CP-element group 695: successors 
    -- CP-element group 695: 	696 
    -- CP-element group 695:  members (5) 
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/word_access_complete/word_0/$exit
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/$exit
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/word_access_complete/word_0/ca
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_Update/word_access_complete/$exit
      -- CP-element group 695: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/ptr_deref_4574_update_completed_
      -- 
    ca_10194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 695_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4574_store_0_ack_1, ack => zeropad3D_CP_2152_elements(695)); -- 
    -- CP-element group 696:  join  transition  place  bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	681 
    -- CP-element group 696: 	689 
    -- CP-element group 696: 	695 
    -- CP-element group 696: successors 
    -- CP-element group 696: 	1120 
    -- CP-element group 696:  members (5) 
      -- CP-element group 696: 	 branch_block_stmt_714/ifx_xelse1397_ifx_xend1445
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576__exit__
      -- CP-element group 696: 	 branch_block_stmt_714/assign_stmt_4476_to_assign_stmt_4576/$exit
      -- CP-element group 696: 	 branch_block_stmt_714/ifx_xelse1397_ifx_xend1445_PhiReq/$exit
      -- CP-element group 696: 	 branch_block_stmt_714/ifx_xelse1397_ifx_xend1445_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_696: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_696"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(681) & zeropad3D_CP_2152_elements(689) & zeropad3D_CP_2152_elements(695);
      gj_zeropad3D_cp_element_group_696 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(696), clk => clk, reset => reset); --
    end block;
    -- CP-element group 697:  transition  input  bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	1120 
    -- CP-element group 697: successors 
    -- CP-element group 697:  members (3) 
      -- CP-element group 697: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Sample/$exit
      -- CP-element group 697: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_sample_completed_
      -- CP-element group 697: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Sample/ra
      -- 
    ra_10206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 697_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4582_inst_ack_0, ack => zeropad3D_CP_2152_elements(697)); -- 
    -- CP-element group 698:  branch  transition  place  input  output  bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	1120 
    -- CP-element group 698: successors 
    -- CP-element group 698: 	699 
    -- CP-element group 698: 	700 
    -- CP-element group 698:  members (13) 
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596__exit__
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597__entry__
      -- CP-element group 698: 	 branch_block_stmt_714/R_cmp1453_4598_place
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_update_completed_
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/$exit
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Update/$exit
      -- CP-element group 698: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Update/ca
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597_dead_link/$entry
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597_eval_test/$entry
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597_eval_test/$exit
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597_eval_test/branch_req
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597_if_link/$entry
      -- CP-element group 698: 	 branch_block_stmt_714/if_stmt_4597_else_link/$entry
      -- 
    ca_10211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4582_inst_ack_1, ack => zeropad3D_CP_2152_elements(698)); -- 
    branch_req_10219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(698), ack => if_stmt_4597_branch_req_0); -- 
    -- CP-element group 699:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	698 
    -- CP-element group 699: successors 
    -- CP-element group 699: 	1129 
    -- CP-element group 699: 	1130 
    -- CP-element group 699: 	1132 
    -- CP-element group 699: 	1133 
    -- CP-element group 699: 	1135 
    -- CP-element group 699: 	1136 
    -- CP-element group 699:  members (40) 
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4609__exit__
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4609__entry__
      -- CP-element group 699: 	 branch_block_stmt_714/merge_stmt_4603__exit__
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xend1445_ifx_xthen1455
      -- CP-element group 699: 	 branch_block_stmt_714/if_stmt_4597_if_link/$exit
      -- CP-element group 699: 	 branch_block_stmt_714/if_stmt_4597_if_link/if_choice_transition
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4609/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/assign_stmt_4609/$exit
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Update/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/merge_stmt_4603_PhiAck/dummy
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/merge_stmt_4603_PhiAck/$exit
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/merge_stmt_4603_PhiAck/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/merge_stmt_4603_PhiReqMerge
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Update/cr
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xend1445_ifx_xthen1455_PhiReq/$exit
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xend1445_ifx_xthen1455_PhiReq/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Update/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Sample/rr
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Sample/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Sample/rr
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Sample/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Update/cr
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Sample/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Sample/rr
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Update/$entry
      -- CP-element group 699: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Update/cr
      -- 
    if_choice_transition_10224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 699_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4597_branch_ack_1, ack => zeropad3D_CP_2152_elements(699)); -- 
    cr_14005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(699), ack => type_cast_4707_inst_req_1); -- 
    rr_14000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(699), ack => type_cast_4707_inst_req_0); -- 
    rr_14023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(699), ack => type_cast_4701_inst_req_0); -- 
    cr_14028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(699), ack => type_cast_4701_inst_req_1); -- 
    rr_14046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(699), ack => type_cast_4694_inst_req_0); -- 
    cr_14051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(699), ack => type_cast_4694_inst_req_1); -- 
    -- CP-element group 700:  fork  transition  place  input  output  bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	698 
    -- CP-element group 700: successors 
    -- CP-element group 700: 	701 
    -- CP-element group 700: 	702 
    -- CP-element group 700: 	703 
    -- CP-element group 700: 	704 
    -- CP-element group 700: 	706 
    -- CP-element group 700: 	709 
    -- CP-element group 700: 	711 
    -- CP-element group 700: 	712 
    -- CP-element group 700: 	713 
    -- CP-element group 700: 	715 
    -- CP-element group 700:  members (54) 
      -- CP-element group 700: 	 branch_block_stmt_714/merge_stmt_4611__exit__
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683__entry__
      -- CP-element group 700: 	 branch_block_stmt_714/merge_stmt_4611_PhiAck/$exit
      -- CP-element group 700: 	 branch_block_stmt_714/ifx_xend1445_ifx_xelse1460
      -- CP-element group 700: 	 branch_block_stmt_714/if_stmt_4597_else_link/$exit
      -- CP-element group 700: 	 branch_block_stmt_714/if_stmt_4597_else_link/else_choice_transition
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_sample_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Sample/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Sample/rr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Update/cr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_sample_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_word_address_calculated
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_root_address_calculated
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/word_access_start/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/word_access_start/word_0/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/word_access_start/word_0/rr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/word_access_complete/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/word_access_complete/word_0/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/word_access_complete/word_0/cr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Update/cr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Update/cr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Update/cr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_sample_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_word_address_calculated
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_root_address_calculated
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/word_access_start/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/word_access_start/word_0/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/word_access_start/word_0/rr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/word_access_complete/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/word_access_complete/word_0/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/word_access_complete/word_0/cr
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_update_start_
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Update/cr
      -- CP-element group 700: 	 branch_block_stmt_714/merge_stmt_4611_PhiAck/dummy
      -- CP-element group 700: 	 branch_block_stmt_714/merge_stmt_4611_PhiAck/$entry
      -- CP-element group 700: 	 branch_block_stmt_714/merge_stmt_4611_PhiReqMerge
      -- CP-element group 700: 	 branch_block_stmt_714/ifx_xend1445_ifx_xelse1460_PhiReq/$exit
      -- CP-element group 700: 	 branch_block_stmt_714/ifx_xend1445_ifx_xelse1460_PhiReq/$entry
      -- 
    else_choice_transition_10228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 700_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4597_branch_ack_0, ack => zeropad3D_CP_2152_elements(700)); -- 
    rr_10244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => type_cast_4621_inst_req_0); -- 
    cr_10249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => type_cast_4621_inst_req_1); -- 
    rr_10266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => LOAD_col_high_4624_load_0_req_0); -- 
    cr_10277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => LOAD_col_high_4624_load_0_req_1); -- 
    cr_10296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => type_cast_4628_inst_req_1); -- 
    cr_10310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => type_cast_4648_inst_req_1); -- 
    cr_10324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => type_cast_4665_inst_req_1); -- 
    rr_10341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => LOAD_row_high_4668_load_0_req_0); -- 
    cr_10352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => LOAD_row_high_4668_load_0_req_1); -- 
    cr_10371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(700), ack => type_cast_4672_inst_req_1); -- 
    -- CP-element group 701:  transition  input  bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	700 
    -- CP-element group 701: successors 
    -- CP-element group 701:  members (3) 
      -- CP-element group 701: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_sample_completed_
      -- CP-element group 701: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Sample/$exit
      -- CP-element group 701: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Sample/ra
      -- 
    ra_10245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 701_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4621_inst_ack_0, ack => zeropad3D_CP_2152_elements(701)); -- 
    -- CP-element group 702:  transition  input  bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	700 
    -- CP-element group 702: successors 
    -- CP-element group 702: 	707 
    -- CP-element group 702:  members (3) 
      -- CP-element group 702: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_update_completed_
      -- CP-element group 702: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Update/$exit
      -- CP-element group 702: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4621_Update/ca
      -- 
    ca_10250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 702_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4621_inst_ack_1, ack => zeropad3D_CP_2152_elements(702)); -- 
    -- CP-element group 703:  transition  input  bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	700 
    -- CP-element group 703: successors 
    -- CP-element group 703:  members (5) 
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_sample_completed_
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/$exit
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/word_access_start/$exit
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/word_access_start/word_0/$exit
      -- CP-element group 703: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Sample/word_access_start/word_0/ra
      -- 
    ra_10267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 703_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4624_load_0_ack_0, ack => zeropad3D_CP_2152_elements(703)); -- 
    -- CP-element group 704:  transition  input  output  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	700 
    -- CP-element group 704: successors 
    -- CP-element group 704: 	705 
    -- CP-element group 704:  members (12) 
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_update_completed_
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/$exit
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/word_access_complete/$exit
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/word_access_complete/word_0/$exit
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/word_access_complete/word_0/ca
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/LOAD_col_high_4624_Merge/$entry
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/LOAD_col_high_4624_Merge/$exit
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/LOAD_col_high_4624_Merge/merge_req
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_col_high_4624_Update/LOAD_col_high_4624_Merge/merge_ack
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_sample_start_
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Sample/$entry
      -- CP-element group 704: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Sample/rr
      -- 
    ca_10278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 704_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4624_load_0_ack_1, ack => zeropad3D_CP_2152_elements(704)); -- 
    rr_10291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(704), ack => type_cast_4628_inst_req_0); -- 
    -- CP-element group 705:  transition  input  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	704 
    -- CP-element group 705: successors 
    -- CP-element group 705:  members (3) 
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_sample_completed_
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Sample/$exit
      -- CP-element group 705: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Sample/ra
      -- 
    ra_10292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 705_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4628_inst_ack_0, ack => zeropad3D_CP_2152_elements(705)); -- 
    -- CP-element group 706:  transition  input  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	700 
    -- CP-element group 706: successors 
    -- CP-element group 706: 	707 
    -- CP-element group 706:  members (3) 
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_update_completed_
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Update/$exit
      -- CP-element group 706: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4628_Update/ca
      -- 
    ca_10297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 706_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4628_inst_ack_1, ack => zeropad3D_CP_2152_elements(706)); -- 
    -- CP-element group 707:  join  transition  output  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	702 
    -- CP-element group 707: 	706 
    -- CP-element group 707: successors 
    -- CP-element group 707: 	708 
    -- CP-element group 707:  members (3) 
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_sample_start_
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Sample/$entry
      -- CP-element group 707: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Sample/rr
      -- 
    rr_10305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(707), ack => type_cast_4648_inst_req_0); -- 
    zeropad3D_cp_element_group_707: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_707"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(702) & zeropad3D_CP_2152_elements(706);
      gj_zeropad3D_cp_element_group_707 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(707), clk => clk, reset => reset); --
    end block;
    -- CP-element group 708:  transition  input  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	707 
    -- CP-element group 708: successors 
    -- CP-element group 708:  members (3) 
      -- CP-element group 708: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_sample_completed_
      -- CP-element group 708: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Sample/$exit
      -- CP-element group 708: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Sample/ra
      -- 
    ra_10306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 708_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4648_inst_ack_0, ack => zeropad3D_CP_2152_elements(708)); -- 
    -- CP-element group 709:  transition  input  output  bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	700 
    -- CP-element group 709: successors 
    -- CP-element group 709: 	710 
    -- CP-element group 709:  members (6) 
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_update_completed_
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Update/$exit
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4648_Update/ca
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_sample_start_
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Sample/$entry
      -- CP-element group 709: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Sample/rr
      -- 
    ca_10311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4648_inst_ack_1, ack => zeropad3D_CP_2152_elements(709)); -- 
    rr_10319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(709), ack => type_cast_4665_inst_req_0); -- 
    -- CP-element group 710:  transition  input  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	709 
    -- CP-element group 710: successors 
    -- CP-element group 710:  members (3) 
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_sample_completed_
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Sample/$exit
      -- CP-element group 710: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Sample/ra
      -- 
    ra_10320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 710_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4665_inst_ack_0, ack => zeropad3D_CP_2152_elements(710)); -- 
    -- CP-element group 711:  transition  input  bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	700 
    -- CP-element group 711: successors 
    -- CP-element group 711: 	716 
    -- CP-element group 711:  members (3) 
      -- CP-element group 711: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_update_completed_
      -- CP-element group 711: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Update/$exit
      -- CP-element group 711: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4665_Update/ca
      -- 
    ca_10325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 711_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4665_inst_ack_1, ack => zeropad3D_CP_2152_elements(711)); -- 
    -- CP-element group 712:  transition  input  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	700 
    -- CP-element group 712: successors 
    -- CP-element group 712:  members (5) 
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_sample_completed_
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/$exit
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/word_access_start/$exit
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/word_access_start/word_0/$exit
      -- CP-element group 712: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Sample/word_access_start/word_0/ra
      -- 
    ra_10342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 712_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4668_load_0_ack_0, ack => zeropad3D_CP_2152_elements(712)); -- 
    -- CP-element group 713:  transition  input  output  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	700 
    -- CP-element group 713: successors 
    -- CP-element group 713: 	714 
    -- CP-element group 713:  members (12) 
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_update_completed_
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/word_access_complete/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/word_access_complete/word_0/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/word_access_complete/word_0/ca
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/LOAD_row_high_4668_Merge/$entry
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/LOAD_row_high_4668_Merge/$exit
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/LOAD_row_high_4668_Merge/merge_req
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/LOAD_row_high_4668_Update/LOAD_row_high_4668_Merge/merge_ack
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_sample_start_
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Sample/$entry
      -- CP-element group 713: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Sample/rr
      -- 
    ca_10353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 713_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4668_load_0_ack_1, ack => zeropad3D_CP_2152_elements(713)); -- 
    rr_10366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(713), ack => type_cast_4672_inst_req_0); -- 
    -- CP-element group 714:  transition  input  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	713 
    -- CP-element group 714: successors 
    -- CP-element group 714:  members (3) 
      -- CP-element group 714: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_sample_completed_
      -- CP-element group 714: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Sample/$exit
      -- CP-element group 714: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Sample/ra
      -- 
    ra_10367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 714_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4672_inst_ack_0, ack => zeropad3D_CP_2152_elements(714)); -- 
    -- CP-element group 715:  transition  input  bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	700 
    -- CP-element group 715: successors 
    -- CP-element group 715: 	716 
    -- CP-element group 715:  members (3) 
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_update_completed_
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Update/$exit
      -- CP-element group 715: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/type_cast_4672_Update/ca
      -- 
    ca_10372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 715_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4672_inst_ack_1, ack => zeropad3D_CP_2152_elements(715)); -- 
    -- CP-element group 716:  branch  join  transition  place  output  bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	711 
    -- CP-element group 716: 	715 
    -- CP-element group 716: successors 
    -- CP-element group 716: 	717 
    -- CP-element group 716: 	718 
    -- CP-element group 716:  members (10) 
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684__entry__
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683__exit__
      -- CP-element group 716: 	 branch_block_stmt_714/R_cmp1487_4685_place
      -- CP-element group 716: 	 branch_block_stmt_714/assign_stmt_4617_to_assign_stmt_4683/$exit
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684_dead_link/$entry
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684_eval_test/$entry
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684_eval_test/$exit
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684_eval_test/branch_req
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684_if_link/$entry
      -- CP-element group 716: 	 branch_block_stmt_714/if_stmt_4684_else_link/$entry
      -- 
    branch_req_10380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(716), ack => if_stmt_4684_branch_req_0); -- 
    zeropad3D_cp_element_group_716: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_716"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(711) & zeropad3D_CP_2152_elements(715);
      gj_zeropad3D_cp_element_group_716 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(716), clk => clk, reset => reset); --
    end block;
    -- CP-element group 717:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	716 
    -- CP-element group 717: successors 
    -- CP-element group 717: 	719 
    -- CP-element group 717: 	720 
    -- CP-element group 717: 	722 
    -- CP-element group 717: 	723 
    -- CP-element group 717: 	724 
    -- CP-element group 717: 	726 
    -- CP-element group 717: 	727 
    -- CP-element group 717: 	728 
    -- CP-element group 717: 	729 
    -- CP-element group 717: 	730 
    -- CP-element group 717: 	731 
    -- CP-element group 717: 	732 
    -- CP-element group 717: 	733 
    -- CP-element group 717: 	734 
    -- CP-element group 717: 	736 
    -- CP-element group 717: 	738 
    -- CP-element group 717: 	740 
    -- CP-element group 717:  members (127) 
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863__entry__
      -- CP-element group 717: 	 branch_block_stmt_714/merge_stmt_4712__exit__
      -- CP-element group 717: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497
      -- CP-element group 717: 	 branch_block_stmt_714/if_stmt_4684_if_link/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/if_stmt_4684_if_link/if_choice_transition
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_word_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_root_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/word_access_start/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/word_access_start/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/word_access_start/word_0/rr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/word_access_complete/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/word_access_complete/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/word_access_complete/word_0/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Update/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_word_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_root_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/word_access_start/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/word_access_start/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/word_access_start/word_0/rr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/word_access_complete/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/word_access_complete/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/word_access_complete/word_0/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Update/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_word_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_root_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/word_access_start/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/word_access_start/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/word_access_start/word_0/rr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/word_access_complete/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/word_access_complete/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/word_access_complete/word_0/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_word_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_root_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/word_access_start/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/word_access_start/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/word_access_start/word_0/rr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/word_access_complete/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/word_access_complete/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/word_access_complete/word_0/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_word_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_root_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_address_resized
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_addr_resize/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_addr_resize/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_addr_resize/base_resize_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_addr_resize/base_resize_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_plus_offset/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_plus_offset/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_plus_offset/sum_rename_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_base_plus_offset/sum_rename_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_word_addrgen/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_word_addrgen/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_word_addrgen/root_register_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_word_addrgen/root_register_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/word_access_start/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/word_access_start/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/word_access_start/word_0/rr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/word_access_complete/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/word_access_complete/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/word_access_complete/word_0/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_sample_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_word_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_root_address_calculated
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_address_resized
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_addr_resize/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_addr_resize/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_addr_resize/base_resize_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_addr_resize/base_resize_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_plus_offset/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_plus_offset/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_plus_offset/sum_rename_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_base_plus_offset/sum_rename_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_word_addrgen/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_word_addrgen/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_word_addrgen/root_register_req
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_word_addrgen/root_register_ack
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/word_access_start/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/word_access_start/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/word_access_start/word_0/rr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/word_access_complete/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/word_access_complete/word_0/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/word_access_complete/word_0/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Update/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Update/cr
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_update_start_
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Update/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Update/cr
      -- CP-element group 717: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/ifx_xelse1460_whilex_xend1497_PhiReq/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/merge_stmt_4712_PhiReqMerge
      -- CP-element group 717: 	 branch_block_stmt_714/merge_stmt_4712_PhiAck/$entry
      -- CP-element group 717: 	 branch_block_stmt_714/merge_stmt_4712_PhiAck/$exit
      -- CP-element group 717: 	 branch_block_stmt_714/merge_stmt_4712_PhiAck/dummy
      -- 
    if_choice_transition_10385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 717_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4684_branch_ack_1, ack => zeropad3D_CP_2152_elements(717)); -- 
    rr_10410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_col_high_4715_load_0_req_0); -- 
    cr_10421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_col_high_4715_load_0_req_1); -- 
    cr_10440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => type_cast_4719_inst_req_1); -- 
    rr_10457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_row_high_4728_load_0_req_0); -- 
    cr_10468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_row_high_4728_load_0_req_1); -- 
    cr_10487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => type_cast_4732_inst_req_1); -- 
    rr_10504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_pad_4747_load_0_req_0); -- 
    cr_10515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_pad_4747_load_0_req_1); -- 
    rr_10537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_depth_high_4750_load_0_req_0); -- 
    cr_10548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => LOAD_depth_high_4750_load_0_req_1); -- 
    rr_10587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => ptr_deref_4762_load_0_req_0); -- 
    cr_10598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => ptr_deref_4762_load_0_req_1); -- 
    rr_10637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => ptr_deref_4774_load_0_req_0); -- 
    cr_10648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => ptr_deref_4774_load_0_req_1); -- 
    cr_10667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => type_cast_4778_inst_req_1); -- 
    cr_10681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => type_cast_4782_inst_req_1); -- 
    cr_10695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(717), ack => type_cast_4821_inst_req_1); -- 
    -- CP-element group 718:  fork  transition  place  input  output  bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	716 
    -- CP-element group 718: successors 
    -- CP-element group 718: 	1121 
    -- CP-element group 718: 	1122 
    -- CP-element group 718: 	1124 
    -- CP-element group 718: 	1125 
    -- CP-element group 718: 	1127 
    -- CP-element group 718:  members (22) 
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496
      -- CP-element group 718: 	 branch_block_stmt_714/if_stmt_4684_else_link/$exit
      -- CP-element group 718: 	 branch_block_stmt_714/if_stmt_4684_else_link/else_choice_transition
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4691/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Update/cr
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Update/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Update/cr
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Update/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Sample/rr
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Sample/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Sample/rr
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/$entry
      -- CP-element group 718: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_10389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 718_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4684_branch_ack_0, ack => zeropad3D_CP_2152_elements(718)); -- 
    cr_13948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(718), ack => type_cast_4709_inst_req_1); -- 
    cr_13971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_13971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(718), ack => type_cast_4703_inst_req_1); -- 
    rr_13966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(718), ack => type_cast_4703_inst_req_0); -- 
    rr_13943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_13943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(718), ack => type_cast_4709_inst_req_0); -- 
    -- CP-element group 719:  transition  input  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	717 
    -- CP-element group 719: successors 
    -- CP-element group 719:  members (5) 
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_sample_completed_
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/$exit
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/word_access_start/$exit
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/word_access_start/word_0/$exit
      -- CP-element group 719: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Sample/word_access_start/word_0/ra
      -- 
    ra_10411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 719_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4715_load_0_ack_0, ack => zeropad3D_CP_2152_elements(719)); -- 
    -- CP-element group 720:  fork  transition  input  output  bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	717 
    -- CP-element group 720: successors 
    -- CP-element group 720: 	721 
    -- CP-element group 720: 	737 
    -- CP-element group 720:  members (15) 
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_update_completed_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/word_access_complete/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/word_access_complete/word_0/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/word_access_complete/word_0/ca
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/LOAD_col_high_4715_Merge/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/LOAD_col_high_4715_Merge/$exit
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/LOAD_col_high_4715_Merge/merge_req
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_col_high_4715_Update/LOAD_col_high_4715_Merge/merge_ack
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_sample_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Sample/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Sample/rr
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_sample_start_
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Sample/$entry
      -- CP-element group 720: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Sample/rr
      -- 
    ca_10422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 720_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4715_load_0_ack_1, ack => zeropad3D_CP_2152_elements(720)); -- 
    rr_10435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => type_cast_4719_inst_req_0); -- 
    rr_10676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(720), ack => type_cast_4782_inst_req_0); -- 
    -- CP-element group 721:  transition  input  bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	720 
    -- CP-element group 721: successors 
    -- CP-element group 721:  members (3) 
      -- CP-element group 721: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_sample_completed_
      -- CP-element group 721: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Sample/$exit
      -- CP-element group 721: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Sample/ra
      -- 
    ra_10436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 721_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4719_inst_ack_0, ack => zeropad3D_CP_2152_elements(721)); -- 
    -- CP-element group 722:  transition  input  bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	717 
    -- CP-element group 722: successors 
    -- CP-element group 722: 	741 
    -- CP-element group 722:  members (3) 
      -- CP-element group 722: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_update_completed_
      -- CP-element group 722: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Update/$exit
      -- CP-element group 722: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4719_Update/ca
      -- 
    ca_10441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4719_inst_ack_1, ack => zeropad3D_CP_2152_elements(722)); -- 
    -- CP-element group 723:  transition  input  bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	717 
    -- CP-element group 723: successors 
    -- CP-element group 723:  members (5) 
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_sample_completed_
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/$exit
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/word_access_start/$exit
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/word_access_start/word_0/$exit
      -- CP-element group 723: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Sample/word_access_start/word_0/ra
      -- 
    ra_10458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 723_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4728_load_0_ack_0, ack => zeropad3D_CP_2152_elements(723)); -- 
    -- CP-element group 724:  transition  input  output  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	717 
    -- CP-element group 724: successors 
    -- CP-element group 724: 	725 
    -- CP-element group 724:  members (12) 
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_update_completed_
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/$exit
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/word_access_complete/$exit
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/word_access_complete/word_0/$exit
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/word_access_complete/word_0/ca
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/LOAD_row_high_4728_Merge/$entry
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/LOAD_row_high_4728_Merge/$exit
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/LOAD_row_high_4728_Merge/merge_req
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_row_high_4728_Update/LOAD_row_high_4728_Merge/merge_ack
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_sample_start_
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Sample/$entry
      -- CP-element group 724: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Sample/rr
      -- 
    ca_10469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 724_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4728_load_0_ack_1, ack => zeropad3D_CP_2152_elements(724)); -- 
    rr_10482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(724), ack => type_cast_4732_inst_req_0); -- 
    -- CP-element group 725:  transition  input  bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	724 
    -- CP-element group 725: successors 
    -- CP-element group 725:  members (3) 
      -- CP-element group 725: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_sample_completed_
      -- CP-element group 725: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Sample/$exit
      -- CP-element group 725: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Sample/ra
      -- 
    ra_10483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4732_inst_ack_0, ack => zeropad3D_CP_2152_elements(725)); -- 
    -- CP-element group 726:  transition  input  bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	717 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	741 
    -- CP-element group 726:  members (3) 
      -- CP-element group 726: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_update_completed_
      -- CP-element group 726: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Update/$exit
      -- CP-element group 726: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4732_Update/ca
      -- 
    ca_10488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 726_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4732_inst_ack_1, ack => zeropad3D_CP_2152_elements(726)); -- 
    -- CP-element group 727:  transition  input  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	717 
    -- CP-element group 727: successors 
    -- CP-element group 727:  members (5) 
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_sample_completed_
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/$exit
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/word_access_start/$exit
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/word_access_start/word_0/$exit
      -- CP-element group 727: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Sample/word_access_start/word_0/ra
      -- 
    ra_10505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 727_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4747_load_0_ack_0, ack => zeropad3D_CP_2152_elements(727)); -- 
    -- CP-element group 728:  transition  input  output  bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	717 
    -- CP-element group 728: successors 
    -- CP-element group 728: 	739 
    -- CP-element group 728:  members (12) 
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_update_completed_
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/word_access_complete/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/word_access_complete/word_0/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/word_access_complete/word_0/ca
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/LOAD_pad_4747_Merge/$entry
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/LOAD_pad_4747_Merge/$exit
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/LOAD_pad_4747_Merge/merge_req
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_pad_4747_Update/LOAD_pad_4747_Merge/merge_ack
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_sample_start_
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Sample/$entry
      -- CP-element group 728: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Sample/rr
      -- 
    ca_10516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_4747_load_0_ack_1, ack => zeropad3D_CP_2152_elements(728)); -- 
    rr_10690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(728), ack => type_cast_4821_inst_req_0); -- 
    -- CP-element group 729:  transition  input  bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	717 
    -- CP-element group 729: successors 
    -- CP-element group 729:  members (5) 
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_sample_completed_
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/$exit
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/word_access_start/$exit
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/word_access_start/word_0/$exit
      -- CP-element group 729: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Sample/word_access_start/word_0/ra
      -- 
    ra_10538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 729_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4750_load_0_ack_0, ack => zeropad3D_CP_2152_elements(729)); -- 
    -- CP-element group 730:  transition  input  output  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	717 
    -- CP-element group 730: successors 
    -- CP-element group 730: 	735 
    -- CP-element group 730:  members (12) 
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_update_completed_
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/$exit
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/word_access_complete/$exit
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/word_access_complete/word_0/$exit
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/word_access_complete/word_0/ca
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/LOAD_depth_high_4750_Merge/$entry
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/LOAD_depth_high_4750_Merge/$exit
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/LOAD_depth_high_4750_Merge/merge_req
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/LOAD_depth_high_4750_Update/LOAD_depth_high_4750_Merge/merge_ack
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_sample_start_
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Sample/$entry
      -- CP-element group 730: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Sample/rr
      -- 
    ca_10549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 730_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_depth_high_4750_load_0_ack_1, ack => zeropad3D_CP_2152_elements(730)); -- 
    rr_10662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(730), ack => type_cast_4778_inst_req_0); -- 
    -- CP-element group 731:  transition  input  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	717 
    -- CP-element group 731: successors 
    -- CP-element group 731:  members (5) 
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_sample_completed_
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/$exit
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/word_access_start/$exit
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/word_access_start/word_0/$exit
      -- CP-element group 731: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Sample/word_access_start/word_0/ra
      -- 
    ra_10588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 731_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4762_load_0_ack_0, ack => zeropad3D_CP_2152_elements(731)); -- 
    -- CP-element group 732:  transition  input  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	717 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	741 
    -- CP-element group 732:  members (9) 
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_update_completed_
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/word_access_complete/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/word_access_complete/word_0/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/word_access_complete/word_0/ca
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/ptr_deref_4762_Merge/$entry
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/ptr_deref_4762_Merge/$exit
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/ptr_deref_4762_Merge/merge_req
      -- CP-element group 732: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4762_Update/ptr_deref_4762_Merge/merge_ack
      -- 
    ca_10599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 732_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4762_load_0_ack_1, ack => zeropad3D_CP_2152_elements(732)); -- 
    -- CP-element group 733:  transition  input  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	717 
    -- CP-element group 733: successors 
    -- CP-element group 733:  members (5) 
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_sample_completed_
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/$exit
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/word_access_start/$exit
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/word_access_start/word_0/$exit
      -- CP-element group 733: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Sample/word_access_start/word_0/ra
      -- 
    ra_10638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 733_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4774_load_0_ack_0, ack => zeropad3D_CP_2152_elements(733)); -- 
    -- CP-element group 734:  transition  input  bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	717 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	741 
    -- CP-element group 734:  members (9) 
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_update_completed_
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/word_access_complete/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/word_access_complete/word_0/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/word_access_complete/word_0/ca
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/ptr_deref_4774_Merge/$entry
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/ptr_deref_4774_Merge/$exit
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/ptr_deref_4774_Merge/merge_req
      -- CP-element group 734: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/ptr_deref_4774_Update/ptr_deref_4774_Merge/merge_ack
      -- 
    ca_10649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 734_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_4774_load_0_ack_1, ack => zeropad3D_CP_2152_elements(734)); -- 
    -- CP-element group 735:  transition  input  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	730 
    -- CP-element group 735: successors 
    -- CP-element group 735:  members (3) 
      -- CP-element group 735: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_sample_completed_
      -- CP-element group 735: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Sample/$exit
      -- CP-element group 735: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Sample/ra
      -- 
    ra_10663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 735_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4778_inst_ack_0, ack => zeropad3D_CP_2152_elements(735)); -- 
    -- CP-element group 736:  transition  input  bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	717 
    -- CP-element group 736: successors 
    -- CP-element group 736: 	741 
    -- CP-element group 736:  members (3) 
      -- CP-element group 736: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_update_completed_
      -- CP-element group 736: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Update/$exit
      -- CP-element group 736: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4778_Update/ca
      -- 
    ca_10668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 736_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4778_inst_ack_1, ack => zeropad3D_CP_2152_elements(736)); -- 
    -- CP-element group 737:  transition  input  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	720 
    -- CP-element group 737: successors 
    -- CP-element group 737:  members (3) 
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_sample_completed_
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Sample/$exit
      -- CP-element group 737: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Sample/ra
      -- 
    ra_10677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 737_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4782_inst_ack_0, ack => zeropad3D_CP_2152_elements(737)); -- 
    -- CP-element group 738:  transition  input  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	717 
    -- CP-element group 738: successors 
    -- CP-element group 738: 	741 
    -- CP-element group 738:  members (3) 
      -- CP-element group 738: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_update_completed_
      -- CP-element group 738: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Update/$exit
      -- CP-element group 738: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4782_Update/ca
      -- 
    ca_10682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 738_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4782_inst_ack_1, ack => zeropad3D_CP_2152_elements(738)); -- 
    -- CP-element group 739:  transition  input  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	728 
    -- CP-element group 739: successors 
    -- CP-element group 739:  members (3) 
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_sample_completed_
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Sample/$exit
      -- CP-element group 739: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Sample/ra
      -- 
    ra_10691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 739_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4821_inst_ack_0, ack => zeropad3D_CP_2152_elements(739)); -- 
    -- CP-element group 740:  transition  input  bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	717 
    -- CP-element group 740: successors 
    -- CP-element group 740: 	741 
    -- CP-element group 740:  members (3) 
      -- CP-element group 740: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_update_completed_
      -- CP-element group 740: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Update/$exit
      -- CP-element group 740: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/type_cast_4821_Update/ca
      -- 
    ca_10696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 740_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4821_inst_ack_1, ack => zeropad3D_CP_2152_elements(740)); -- 
    -- CP-element group 741:  join  fork  transition  place  output  bypass 
    -- CP-element group 741: predecessors 
    -- CP-element group 741: 	722 
    -- CP-element group 741: 	726 
    -- CP-element group 741: 	732 
    -- CP-element group 741: 	734 
    -- CP-element group 741: 	736 
    -- CP-element group 741: 	738 
    -- CP-element group 741: 	740 
    -- CP-element group 741: successors 
    -- CP-element group 741: 	1154 
    -- CP-element group 741: 	1155 
    -- CP-element group 741: 	1157 
    -- CP-element group 741: 	1158 
    -- CP-element group 741: 	1160 
    -- CP-element group 741:  members (22) 
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863__exit__
      -- CP-element group 741: 	 branch_block_stmt_714/assign_stmt_4716_to_assign_stmt_4863/$exit
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Sample/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Sample/rr
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Update/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Update/cr
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Sample/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Sample/rr
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Update/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Update/cr
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4866/$entry
      -- CP-element group 741: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/$entry
      -- 
    rr_14159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(741), ack => type_cast_4882_inst_req_0); -- 
    cr_14164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(741), ack => type_cast_4882_inst_req_1); -- 
    rr_14182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(741), ack => type_cast_4878_inst_req_0); -- 
    cr_14187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(741), ack => type_cast_4878_inst_req_1); -- 
    zeropad3D_cp_element_group_741: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_741"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(722) & zeropad3D_CP_2152_elements(726) & zeropad3D_CP_2152_elements(732) & zeropad3D_CP_2152_elements(734) & zeropad3D_CP_2152_elements(736) & zeropad3D_CP_2152_elements(738) & zeropad3D_CP_2152_elements(740);
      gj_zeropad3D_cp_element_group_741 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(741), clk => clk, reset => reset); --
    end block;
    -- CP-element group 742:  transition  input  bypass 
    -- CP-element group 742: predecessors 
    -- CP-element group 742: 	1166 
    -- CP-element group 742: successors 
    -- CP-element group 742:  members (3) 
      -- CP-element group 742: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_sample_completed_
      -- CP-element group 742: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Sample/$exit
      -- CP-element group 742: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Sample/ra
      -- 
    ra_10708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 742_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4889_inst_ack_0, ack => zeropad3D_CP_2152_elements(742)); -- 
    -- CP-element group 743:  branch  transition  place  input  output  bypass 
    -- CP-element group 743: predecessors 
    -- CP-element group 743: 	1166 
    -- CP-element group 743: successors 
    -- CP-element group 743: 	744 
    -- CP-element group 743: 	745 
    -- CP-element group 743:  members (13) 
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897__exit__
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898__entry__
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_update_completed_
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Update/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Update/ca
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898_dead_link/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898_eval_test/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898_eval_test/$exit
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898_eval_test/branch_req
      -- CP-element group 743: 	 branch_block_stmt_714/R_cmp1567_4899_place
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898_if_link/$entry
      -- CP-element group 743: 	 branch_block_stmt_714/if_stmt_4898_else_link/$entry
      -- 
    ca_10713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 743_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4889_inst_ack_1, ack => zeropad3D_CP_2152_elements(743)); -- 
    branch_req_10721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(743), ack => if_stmt_4898_branch_req_0); -- 
    -- CP-element group 744:  transition  place  input  bypass 
    -- CP-element group 744: predecessors 
    -- CP-element group 744: 	743 
    -- CP-element group 744: successors 
    -- CP-element group 744: 	1167 
    -- CP-element group 744:  members (5) 
      -- CP-element group 744: 	 branch_block_stmt_714/if_stmt_4898_if_link/$exit
      -- CP-element group 744: 	 branch_block_stmt_714/if_stmt_4898_if_link/if_choice_transition
      -- CP-element group 744: 	 branch_block_stmt_714/whilex_xbody1562_ifx_xthen1596
      -- CP-element group 744: 	 branch_block_stmt_714/whilex_xbody1562_ifx_xthen1596_PhiReq/$entry
      -- CP-element group 744: 	 branch_block_stmt_714/whilex_xbody1562_ifx_xthen1596_PhiReq/$exit
      -- 
    if_choice_transition_10726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 744_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4898_branch_ack_1, ack => zeropad3D_CP_2152_elements(744)); -- 
    -- CP-element group 745:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 745: predecessors 
    -- CP-element group 745: 	743 
    -- CP-element group 745: successors 
    -- CP-element group 745: 	746 
    -- CP-element group 745: 	747 
    -- CP-element group 745: 	749 
    -- CP-element group 745:  members (27) 
      -- CP-element group 745: 	 branch_block_stmt_714/merge_stmt_4904__exit__
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923__entry__
      -- CP-element group 745: 	 branch_block_stmt_714/if_stmt_4898_else_link/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/if_stmt_4898_else_link/else_choice_transition
      -- CP-element group 745: 	 branch_block_stmt_714/whilex_xbody1562_lorx_xlhsx_xfalse1569
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_sample_start_
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_update_start_
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_word_address_calculated
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_root_address_calculated
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/word_access_start/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/word_access_start/word_0/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/word_access_start/word_0/rr
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/word_access_complete/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/word_access_complete/word_0/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/word_access_complete/word_0/cr
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_update_start_
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Update/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Update/cr
      -- CP-element group 745: 	 branch_block_stmt_714/whilex_xbody1562_lorx_xlhsx_xfalse1569_PhiReq/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/whilex_xbody1562_lorx_xlhsx_xfalse1569_PhiReq/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/merge_stmt_4904_PhiReqMerge
      -- CP-element group 745: 	 branch_block_stmt_714/merge_stmt_4904_PhiAck/$entry
      -- CP-element group 745: 	 branch_block_stmt_714/merge_stmt_4904_PhiAck/$exit
      -- CP-element group 745: 	 branch_block_stmt_714/merge_stmt_4904_PhiAck/dummy
      -- 
    else_choice_transition_10730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 745_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4898_branch_ack_0, ack => zeropad3D_CP_2152_elements(745)); -- 
    rr_10751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(745), ack => LOAD_row_high_4906_load_0_req_0); -- 
    cr_10762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(745), ack => LOAD_row_high_4906_load_0_req_1); -- 
    cr_10781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(745), ack => type_cast_4910_inst_req_1); -- 
    -- CP-element group 746:  transition  input  bypass 
    -- CP-element group 746: predecessors 
    -- CP-element group 746: 	745 
    -- CP-element group 746: successors 
    -- CP-element group 746:  members (5) 
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_sample_completed_
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/$exit
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/word_access_start/$exit
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/word_access_start/word_0/$exit
      -- CP-element group 746: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Sample/word_access_start/word_0/ra
      -- 
    ra_10752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 746_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4906_load_0_ack_0, ack => zeropad3D_CP_2152_elements(746)); -- 
    -- CP-element group 747:  transition  input  output  bypass 
    -- CP-element group 747: predecessors 
    -- CP-element group 747: 	745 
    -- CP-element group 747: successors 
    -- CP-element group 747: 	748 
    -- CP-element group 747:  members (12) 
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_update_completed_
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/word_access_complete/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/word_access_complete/word_0/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/word_access_complete/word_0/ca
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/LOAD_row_high_4906_Merge/$entry
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/LOAD_row_high_4906_Merge/$exit
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/LOAD_row_high_4906_Merge/merge_req
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/LOAD_row_high_4906_Update/LOAD_row_high_4906_Merge/merge_ack
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_sample_start_
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Sample/$entry
      -- CP-element group 747: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Sample/rr
      -- 
    ca_10763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 747_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_4906_load_0_ack_1, ack => zeropad3D_CP_2152_elements(747)); -- 
    rr_10776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(747), ack => type_cast_4910_inst_req_0); -- 
    -- CP-element group 748:  transition  input  bypass 
    -- CP-element group 748: predecessors 
    -- CP-element group 748: 	747 
    -- CP-element group 748: successors 
    -- CP-element group 748:  members (3) 
      -- CP-element group 748: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_sample_completed_
      -- CP-element group 748: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Sample/$exit
      -- CP-element group 748: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Sample/ra
      -- 
    ra_10777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 748_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4910_inst_ack_0, ack => zeropad3D_CP_2152_elements(748)); -- 
    -- CP-element group 749:  branch  transition  place  input  output  bypass 
    -- CP-element group 749: predecessors 
    -- CP-element group 749: 	745 
    -- CP-element group 749: successors 
    -- CP-element group 749: 	750 
    -- CP-element group 749: 	751 
    -- CP-element group 749:  members (13) 
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923__exit__
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924__entry__
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/$exit
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_update_completed_
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Update/$exit
      -- CP-element group 749: 	 branch_block_stmt_714/assign_stmt_4907_to_assign_stmt_4923/type_cast_4910_Update/ca
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924_dead_link/$entry
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924_eval_test/$entry
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924_eval_test/$exit
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924_eval_test/branch_req
      -- CP-element group 749: 	 branch_block_stmt_714/R_cmp1577_4925_place
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924_if_link/$entry
      -- CP-element group 749: 	 branch_block_stmt_714/if_stmt_4924_else_link/$entry
      -- 
    ca_10782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 749_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4910_inst_ack_1, ack => zeropad3D_CP_2152_elements(749)); -- 
    branch_req_10790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(749), ack => if_stmt_4924_branch_req_0); -- 
    -- CP-element group 750:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 750: predecessors 
    -- CP-element group 750: 	749 
    -- CP-element group 750: successors 
    -- CP-element group 750: 	752 
    -- CP-element group 750: 	753 
    -- CP-element group 750:  members (18) 
      -- CP-element group 750: 	 branch_block_stmt_714/merge_stmt_4930__exit__
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942__entry__
      -- CP-element group 750: 	 branch_block_stmt_714/if_stmt_4924_if_link/$exit
      -- CP-element group 750: 	 branch_block_stmt_714/if_stmt_4924_if_link/if_choice_transition
      -- CP-element group 750: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1579
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/$entry
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_sample_start_
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_update_start_
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Sample/$entry
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Sample/rr
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Update/$entry
      -- CP-element group 750: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Update/cr
      -- CP-element group 750: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1579_PhiReq/$entry
      -- CP-element group 750: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_lorx_xlhsx_xfalse1579_PhiReq/$exit
      -- CP-element group 750: 	 branch_block_stmt_714/merge_stmt_4930_PhiReqMerge
      -- CP-element group 750: 	 branch_block_stmt_714/merge_stmt_4930_PhiAck/$entry
      -- CP-element group 750: 	 branch_block_stmt_714/merge_stmt_4930_PhiAck/$exit
      -- CP-element group 750: 	 branch_block_stmt_714/merge_stmt_4930_PhiAck/dummy
      -- 
    if_choice_transition_10795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 750_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4924_branch_ack_1, ack => zeropad3D_CP_2152_elements(750)); -- 
    rr_10812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(750), ack => type_cast_4934_inst_req_0); -- 
    cr_10817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(750), ack => type_cast_4934_inst_req_1); -- 
    -- CP-element group 751:  transition  place  input  bypass 
    -- CP-element group 751: predecessors 
    -- CP-element group 751: 	749 
    -- CP-element group 751: successors 
    -- CP-element group 751: 	1167 
    -- CP-element group 751:  members (5) 
      -- CP-element group 751: 	 branch_block_stmt_714/if_stmt_4924_else_link/$exit
      -- CP-element group 751: 	 branch_block_stmt_714/if_stmt_4924_else_link/else_choice_transition
      -- CP-element group 751: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_ifx_xthen1596
      -- CP-element group 751: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_ifx_xthen1596_PhiReq/$entry
      -- CP-element group 751: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1569_ifx_xthen1596_PhiReq/$exit
      -- 
    else_choice_transition_10799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 751_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4924_branch_ack_0, ack => zeropad3D_CP_2152_elements(751)); -- 
    -- CP-element group 752:  transition  input  bypass 
    -- CP-element group 752: predecessors 
    -- CP-element group 752: 	750 
    -- CP-element group 752: successors 
    -- CP-element group 752:  members (3) 
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_sample_completed_
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Sample/$exit
      -- CP-element group 752: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Sample/ra
      -- 
    ra_10813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 752_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4934_inst_ack_0, ack => zeropad3D_CP_2152_elements(752)); -- 
    -- CP-element group 753:  branch  transition  place  input  output  bypass 
    -- CP-element group 753: predecessors 
    -- CP-element group 753: 	750 
    -- CP-element group 753: successors 
    -- CP-element group 753: 	754 
    -- CP-element group 753: 	755 
    -- CP-element group 753:  members (13) 
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942__exit__
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943__entry__
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/$exit
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_update_completed_
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Update/$exit
      -- CP-element group 753: 	 branch_block_stmt_714/assign_stmt_4935_to_assign_stmt_4942/type_cast_4934_Update/ca
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943_dead_link/$entry
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943_eval_test/$entry
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943_eval_test/$exit
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943_eval_test/branch_req
      -- CP-element group 753: 	 branch_block_stmt_714/R_cmp1584_4944_place
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943_if_link/$entry
      -- CP-element group 753: 	 branch_block_stmt_714/if_stmt_4943_else_link/$entry
      -- 
    ca_10818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 753_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4934_inst_ack_1, ack => zeropad3D_CP_2152_elements(753)); -- 
    branch_req_10826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(753), ack => if_stmt_4943_branch_req_0); -- 
    -- CP-element group 754:  transition  place  input  bypass 
    -- CP-element group 754: predecessors 
    -- CP-element group 754: 	753 
    -- CP-element group 754: successors 
    -- CP-element group 754: 	1167 
    -- CP-element group 754:  members (5) 
      -- CP-element group 754: 	 branch_block_stmt_714/if_stmt_4943_if_link/$exit
      -- CP-element group 754: 	 branch_block_stmt_714/if_stmt_4943_if_link/if_choice_transition
      -- CP-element group 754: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_ifx_xthen1596
      -- CP-element group 754: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_ifx_xthen1596_PhiReq/$entry
      -- CP-element group 754: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_ifx_xthen1596_PhiReq/$exit
      -- 
    if_choice_transition_10831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 754_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4943_branch_ack_1, ack => zeropad3D_CP_2152_elements(754)); -- 
    -- CP-element group 755:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 755: predecessors 
    -- CP-element group 755: 	753 
    -- CP-element group 755: successors 
    -- CP-element group 755: 	756 
    -- CP-element group 755: 	757 
    -- CP-element group 755: 	759 
    -- CP-element group 755:  members (27) 
      -- CP-element group 755: 	 branch_block_stmt_714/merge_stmt_4949__exit__
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968__entry__
      -- CP-element group 755: 	 branch_block_stmt_714/if_stmt_4943_else_link/$exit
      -- CP-element group 755: 	 branch_block_stmt_714/if_stmt_4943_else_link/else_choice_transition
      -- CP-element group 755: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_lorx_xlhsx_xfalse1586
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_sample_start_
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_update_start_
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_word_address_calculated
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_root_address_calculated
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/word_access_start/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/word_access_start/word_0/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/word_access_start/word_0/rr
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/word_access_complete/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/word_access_complete/word_0/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/word_access_complete/word_0/cr
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_update_start_
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Update/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Update/cr
      -- CP-element group 755: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_lorx_xlhsx_xfalse1586_PhiReq/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1579_lorx_xlhsx_xfalse1586_PhiReq/$exit
      -- CP-element group 755: 	 branch_block_stmt_714/merge_stmt_4949_PhiReqMerge
      -- CP-element group 755: 	 branch_block_stmt_714/merge_stmt_4949_PhiAck/$entry
      -- CP-element group 755: 	 branch_block_stmt_714/merge_stmt_4949_PhiAck/$exit
      -- CP-element group 755: 	 branch_block_stmt_714/merge_stmt_4949_PhiAck/dummy
      -- 
    else_choice_transition_10835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 755_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4943_branch_ack_0, ack => zeropad3D_CP_2152_elements(755)); -- 
    rr_10856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(755), ack => LOAD_col_high_4951_load_0_req_0); -- 
    cr_10867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(755), ack => LOAD_col_high_4951_load_0_req_1); -- 
    cr_10886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(755), ack => type_cast_4955_inst_req_1); -- 
    -- CP-element group 756:  transition  input  bypass 
    -- CP-element group 756: predecessors 
    -- CP-element group 756: 	755 
    -- CP-element group 756: successors 
    -- CP-element group 756:  members (5) 
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_sample_completed_
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/$exit
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/word_access_start/$exit
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/word_access_start/word_0/$exit
      -- CP-element group 756: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Sample/word_access_start/word_0/ra
      -- 
    ra_10857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 756_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4951_load_0_ack_0, ack => zeropad3D_CP_2152_elements(756)); -- 
    -- CP-element group 757:  transition  input  output  bypass 
    -- CP-element group 757: predecessors 
    -- CP-element group 757: 	755 
    -- CP-element group 757: successors 
    -- CP-element group 757: 	758 
    -- CP-element group 757:  members (12) 
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_update_completed_
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/word_access_complete/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/word_access_complete/word_0/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/word_access_complete/word_0/ca
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/LOAD_col_high_4951_Merge/$entry
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/LOAD_col_high_4951_Merge/$exit
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/LOAD_col_high_4951_Merge/merge_req
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/LOAD_col_high_4951_Update/LOAD_col_high_4951_Merge/merge_ack
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_sample_start_
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Sample/$entry
      -- CP-element group 757: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Sample/rr
      -- 
    ca_10868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 757_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_4951_load_0_ack_1, ack => zeropad3D_CP_2152_elements(757)); -- 
    rr_10881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(757), ack => type_cast_4955_inst_req_0); -- 
    -- CP-element group 758:  transition  input  bypass 
    -- CP-element group 758: predecessors 
    -- CP-element group 758: 	757 
    -- CP-element group 758: successors 
    -- CP-element group 758:  members (3) 
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_sample_completed_
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Sample/$exit
      -- CP-element group 758: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Sample/ra
      -- 
    ra_10882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 758_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4955_inst_ack_0, ack => zeropad3D_CP_2152_elements(758)); -- 
    -- CP-element group 759:  branch  transition  place  input  output  bypass 
    -- CP-element group 759: predecessors 
    -- CP-element group 759: 	755 
    -- CP-element group 759: successors 
    -- CP-element group 759: 	760 
    -- CP-element group 759: 	761 
    -- CP-element group 759:  members (13) 
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968__exit__
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969__entry__
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969_else_link/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969_if_link/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969_eval_test/branch_req
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969_eval_test/$exit
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969_eval_test/$entry
      -- CP-element group 759: 	 branch_block_stmt_714/R_cmp1594_4970_place
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/$exit
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_update_completed_
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Update/$exit
      -- CP-element group 759: 	 branch_block_stmt_714/assign_stmt_4952_to_assign_stmt_4968/type_cast_4955_Update/ca
      -- CP-element group 759: 	 branch_block_stmt_714/if_stmt_4969_dead_link/$entry
      -- 
    ca_10887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 759_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4955_inst_ack_1, ack => zeropad3D_CP_2152_elements(759)); -- 
    branch_req_10895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_10895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(759), ack => if_stmt_4969_branch_req_0); -- 
    -- CP-element group 760:  fork  transition  place  input  output  bypass 
    -- CP-element group 760: predecessors 
    -- CP-element group 760: 	759 
    -- CP-element group 760: successors 
    -- CP-element group 760: 	776 
    -- CP-element group 760: 	777 
    -- CP-element group 760: 	779 
    -- CP-element group 760: 	781 
    -- CP-element group 760: 	783 
    -- CP-element group 760: 	785 
    -- CP-element group 760: 	787 
    -- CP-element group 760: 	789 
    -- CP-element group 760: 	791 
    -- CP-element group 760: 	794 
    -- CP-element group 760:  members (46) 
      -- CP-element group 760: 	 branch_block_stmt_714/merge_stmt_5033__exit__
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138__entry__
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Sample/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Sample/rr
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/if_stmt_4969_if_link/$exit
      -- CP-element group 760: 	 branch_block_stmt_714/if_stmt_4969_if_link/if_choice_transition
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Update/cr
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/word_access_complete/word_0/cr
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/word_access_complete/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/word_access_complete/word_0/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/word_access_complete/word_0/cr
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Update/req
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Update/cr
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/word_access_complete/word_0/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_sample_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Update/cr
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Update/req
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_update_start
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Update/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_update_start
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_update_start_
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_complete/req
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_complete/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xelse1617
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_complete/req
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/word_access_complete/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_complete/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xelse1617_PhiReq/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xelse1617_PhiReq/$exit
      -- CP-element group 760: 	 branch_block_stmt_714/merge_stmt_5033_PhiReqMerge
      -- CP-element group 760: 	 branch_block_stmt_714/merge_stmt_5033_PhiAck/$entry
      -- CP-element group 760: 	 branch_block_stmt_714/merge_stmt_5033_PhiAck/$exit
      -- CP-element group 760: 	 branch_block_stmt_714/merge_stmt_5033_PhiAck/dummy
      -- 
    if_choice_transition_10900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 760_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4969_branch_ack_1, ack => zeropad3D_CP_2152_elements(760)); -- 
    rr_11058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => type_cast_5037_inst_req_0); -- 
    cr_11063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => type_cast_5037_inst_req_1); -- 
    cr_11283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => ptr_deref_5136_store_0_req_1); -- 
    cr_11168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => ptr_deref_5112_load_0_req_1); -- 
    req_11218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => array_obj_ref_5132_index_offset_req_1); -- 
    cr_11077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => type_cast_5101_inst_req_1); -- 
    cr_11187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => type_cast_5126_inst_req_1); -- 
    req_11108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => array_obj_ref_5107_index_offset_req_1); -- 
    req_11233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => addr_of_5133_final_reg_req_1); -- 
    req_11123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(760), ack => addr_of_5108_final_reg_req_1); -- 
    -- CP-element group 761:  transition  place  input  bypass 
    -- CP-element group 761: predecessors 
    -- CP-element group 761: 	759 
    -- CP-element group 761: successors 
    -- CP-element group 761: 	1167 
    -- CP-element group 761:  members (5) 
      -- CP-element group 761: 	 branch_block_stmt_714/if_stmt_4969_else_link/$exit
      -- CP-element group 761: 	 branch_block_stmt_714/if_stmt_4969_else_link/else_choice_transition
      -- CP-element group 761: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xthen1596
      -- CP-element group 761: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xthen1596_PhiReq/$entry
      -- CP-element group 761: 	 branch_block_stmt_714/lorx_xlhsx_xfalse1586_ifx_xthen1596_PhiReq/$exit
      -- 
    else_choice_transition_10904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 761_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_4969_branch_ack_0, ack => zeropad3D_CP_2152_elements(761)); -- 
    -- CP-element group 762:  transition  input  bypass 
    -- CP-element group 762: predecessors 
    -- CP-element group 762: 	1167 
    -- CP-element group 762: successors 
    -- CP-element group 762:  members (3) 
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_sample_completed_
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Sample/ra
      -- CP-element group 762: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Sample/$exit
      -- 
    ra_10918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 762_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4979_inst_ack_0, ack => zeropad3D_CP_2152_elements(762)); -- 
    -- CP-element group 763:  transition  input  bypass 
    -- CP-element group 763: predecessors 
    -- CP-element group 763: 	1167 
    -- CP-element group 763: successors 
    -- CP-element group 763: 	766 
    -- CP-element group 763:  members (3) 
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_update_completed_
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Update/ca
      -- CP-element group 763: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Update/$exit
      -- 
    ca_10923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 763_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4979_inst_ack_1, ack => zeropad3D_CP_2152_elements(763)); -- 
    -- CP-element group 764:  transition  input  bypass 
    -- CP-element group 764: predecessors 
    -- CP-element group 764: 	1167 
    -- CP-element group 764: successors 
    -- CP-element group 764:  members (3) 
      -- CP-element group 764: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Sample/ra
      -- CP-element group 764: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Sample/$exit
      -- CP-element group 764: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_sample_completed_
      -- 
    ra_10932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 764_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4984_inst_ack_0, ack => zeropad3D_CP_2152_elements(764)); -- 
    -- CP-element group 765:  transition  input  bypass 
    -- CP-element group 765: predecessors 
    -- CP-element group 765: 	1167 
    -- CP-element group 765: successors 
    -- CP-element group 765: 	766 
    -- CP-element group 765:  members (3) 
      -- CP-element group 765: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Update/ca
      -- CP-element group 765: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Update/$exit
      -- CP-element group 765: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_update_completed_
      -- 
    ca_10937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 765_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4984_inst_ack_1, ack => zeropad3D_CP_2152_elements(765)); -- 
    -- CP-element group 766:  join  transition  output  bypass 
    -- CP-element group 766: predecessors 
    -- CP-element group 766: 	763 
    -- CP-element group 766: 	765 
    -- CP-element group 766: successors 
    -- CP-element group 766: 	767 
    -- CP-element group 766:  members (3) 
      -- CP-element group 766: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Sample/rr
      -- CP-element group 766: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Sample/$entry
      -- CP-element group 766: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_sample_start_
      -- 
    rr_10945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(766), ack => type_cast_5018_inst_req_0); -- 
    zeropad3D_cp_element_group_766: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_766"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(763) & zeropad3D_CP_2152_elements(765);
      gj_zeropad3D_cp_element_group_766 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(766), clk => clk, reset => reset); --
    end block;
    -- CP-element group 767:  transition  input  bypass 
    -- CP-element group 767: predecessors 
    -- CP-element group 767: 	766 
    -- CP-element group 767: successors 
    -- CP-element group 767:  members (3) 
      -- CP-element group 767: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Sample/ra
      -- CP-element group 767: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Sample/$exit
      -- CP-element group 767: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_sample_completed_
      -- 
    ra_10946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 767_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5018_inst_ack_0, ack => zeropad3D_CP_2152_elements(767)); -- 
    -- CP-element group 768:  transition  input  output  bypass 
    -- CP-element group 768: predecessors 
    -- CP-element group 768: 	1167 
    -- CP-element group 768: successors 
    -- CP-element group 768: 	769 
    -- CP-element group 768:  members (16) 
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_scale_1/$exit
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_scale_1/scale_rename_req
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_scale_1/scale_rename_ack
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_resized_1
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_scaled_1
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Sample/$entry
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Sample/req
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_computed_1
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_resize_1/$entry
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_resize_1/$exit
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_resize_1/index_resize_req
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_resize_1/index_resize_ack
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Update/ca
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Update/$exit
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_update_completed_
      -- CP-element group 768: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_index_scale_1/$entry
      -- 
    ca_10951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 768_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5018_inst_ack_1, ack => zeropad3D_CP_2152_elements(768)); -- 
    req_10976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(768), ack => array_obj_ref_5024_index_offset_req_0); -- 
    -- CP-element group 769:  transition  input  bypass 
    -- CP-element group 769: predecessors 
    -- CP-element group 769: 	768 
    -- CP-element group 769: successors 
    -- CP-element group 769: 	775 
    -- CP-element group 769:  members (3) 
      -- CP-element group 769: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_sample_complete
      -- CP-element group 769: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Sample/$exit
      -- CP-element group 769: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Sample/ack
      -- 
    ack_10977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 769_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5024_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(769)); -- 
    -- CP-element group 770:  transition  input  output  bypass 
    -- CP-element group 770: predecessors 
    -- CP-element group 770: 	1167 
    -- CP-element group 770: successors 
    -- CP-element group 770: 	771 
    -- CP-element group 770:  members (11) 
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_root_address_calculated
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_offset_calculated
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Update/$exit
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Update/ack
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_base_plus_offset/$entry
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_base_plus_offset/$exit
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_base_plus_offset/sum_rename_req
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_base_plus_offset/sum_rename_ack
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_sample_start_
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_request/req
      -- CP-element group 770: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_request/$entry
      -- 
    ack_10982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 770_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5024_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(770)); -- 
    req_10991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(770), ack => addr_of_5025_final_reg_req_0); -- 
    -- CP-element group 771:  transition  input  bypass 
    -- CP-element group 771: predecessors 
    -- CP-element group 771: 	770 
    -- CP-element group 771: successors 
    -- CP-element group 771:  members (3) 
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_sample_completed_
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_request/ack
      -- CP-element group 771: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_request/$exit
      -- 
    ack_10992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 771_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5025_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(771)); -- 
    -- CP-element group 772:  join  fork  transition  input  output  bypass 
    -- CP-element group 772: predecessors 
    -- CP-element group 772: 	1167 
    -- CP-element group 772: successors 
    -- CP-element group 772: 	773 
    -- CP-element group 772:  members (28) 
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_address_calculated
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_word_address_calculated
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_update_completed_
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_root_address_calculated
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_address_resized
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_addr_resize/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_addr_resize/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_addr_resize/base_resize_req
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_addr_resize/base_resize_ack
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_plus_offset/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_plus_offset/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_plus_offset/sum_rename_req
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_sample_start_
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_complete/ack
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_complete/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/word_access_start/word_0/rr
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/word_access_start/word_0/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/word_access_start/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/ptr_deref_5028_Split/split_ack
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/ptr_deref_5028_Split/split_req
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/ptr_deref_5028_Split/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/ptr_deref_5028_Split/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_word_addrgen/root_register_ack
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_word_addrgen/root_register_req
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_word_addrgen/$exit
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_word_addrgen/$entry
      -- CP-element group 772: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_base_plus_offset/sum_rename_ack
      -- 
    ack_10997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 772_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5025_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(772)); -- 
    rr_11035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(772), ack => ptr_deref_5028_store_0_req_0); -- 
    -- CP-element group 773:  transition  input  bypass 
    -- CP-element group 773: predecessors 
    -- CP-element group 773: 	772 
    -- CP-element group 773: successors 
    -- CP-element group 773:  members (5) 
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_sample_completed_
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/word_access_start/word_0/ra
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/word_access_start/word_0/$exit
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/word_access_start/$exit
      -- CP-element group 773: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Sample/$exit
      -- 
    ra_11036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 773_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5028_store_0_ack_0, ack => zeropad3D_CP_2152_elements(773)); -- 
    -- CP-element group 774:  transition  input  bypass 
    -- CP-element group 774: predecessors 
    -- CP-element group 774: 	1167 
    -- CP-element group 774: successors 
    -- CP-element group 774: 	775 
    -- CP-element group 774:  members (5) 
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_update_completed_
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/word_access_complete/word_0/ca
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/word_access_complete/word_0/$exit
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/word_access_complete/$exit
      -- CP-element group 774: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/$exit
      -- 
    ca_11047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 774_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5028_store_0_ack_1, ack => zeropad3D_CP_2152_elements(774)); -- 
    -- CP-element group 775:  join  transition  place  bypass 
    -- CP-element group 775: predecessors 
    -- CP-element group 775: 	769 
    -- CP-element group 775: 	774 
    -- CP-element group 775: successors 
    -- CP-element group 775: 	1168 
    -- CP-element group 775:  members (5) 
      -- CP-element group 775: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031__exit__
      -- CP-element group 775: 	 branch_block_stmt_714/ifx_xthen1596_ifx_xend1665
      -- CP-element group 775: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/$exit
      -- CP-element group 775: 	 branch_block_stmt_714/ifx_xthen1596_ifx_xend1665_PhiReq/$entry
      -- CP-element group 775: 	 branch_block_stmt_714/ifx_xthen1596_ifx_xend1665_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_775: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_775"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(769) & zeropad3D_CP_2152_elements(774);
      gj_zeropad3D_cp_element_group_775 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(775), clk => clk, reset => reset); --
    end block;
    -- CP-element group 776:  transition  input  bypass 
    -- CP-element group 776: predecessors 
    -- CP-element group 776: 	760 
    -- CP-element group 776: successors 
    -- CP-element group 776:  members (3) 
      -- CP-element group 776: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Sample/$exit
      -- CP-element group 776: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Sample/ra
      -- CP-element group 776: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_sample_completed_
      -- 
    ra_11059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 776_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5037_inst_ack_0, ack => zeropad3D_CP_2152_elements(776)); -- 
    -- CP-element group 777:  fork  transition  input  output  bypass 
    -- CP-element group 777: predecessors 
    -- CP-element group 777: 	760 
    -- CP-element group 777: successors 
    -- CP-element group 777: 	778 
    -- CP-element group 777: 	786 
    -- CP-element group 777:  members (9) 
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Update/$exit
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_Update/ca
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_sample_start_
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Sample/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Sample/rr
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5037_update_completed_
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Sample/rr
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Sample/$entry
      -- CP-element group 777: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_sample_start_
      -- 
    ca_11064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 777_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5037_inst_ack_1, ack => zeropad3D_CP_2152_elements(777)); -- 
    rr_11072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(777), ack => type_cast_5101_inst_req_0); -- 
    rr_11182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(777), ack => type_cast_5126_inst_req_0); -- 
    -- CP-element group 778:  transition  input  bypass 
    -- CP-element group 778: predecessors 
    -- CP-element group 778: 	777 
    -- CP-element group 778: successors 
    -- CP-element group 778:  members (3) 
      -- CP-element group 778: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_sample_completed_
      -- CP-element group 778: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Sample/$exit
      -- CP-element group 778: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Sample/ra
      -- 
    ra_11073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 778_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5101_inst_ack_0, ack => zeropad3D_CP_2152_elements(778)); -- 
    -- CP-element group 779:  transition  input  output  bypass 
    -- CP-element group 779: predecessors 
    -- CP-element group 779: 	760 
    -- CP-element group 779: successors 
    -- CP-element group 779: 	780 
    -- CP-element group 779:  members (16) 
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_update_completed_
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Update/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5101_Update/ca
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Sample/req
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Sample/$entry
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_scale_1/scale_rename_ack
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_scale_1/scale_rename_req
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_scale_1/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_scale_1/$entry
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_resize_1/index_resize_ack
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_resize_1/index_resize_req
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_resize_1/$exit
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_resize_1/$entry
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_computed_1
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_scaled_1
      -- CP-element group 779: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_index_resized_1
      -- 
    ca_11078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 779_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5101_inst_ack_1, ack => zeropad3D_CP_2152_elements(779)); -- 
    req_11103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(779), ack => array_obj_ref_5107_index_offset_req_0); -- 
    -- CP-element group 780:  transition  input  bypass 
    -- CP-element group 780: predecessors 
    -- CP-element group 780: 	779 
    -- CP-element group 780: successors 
    -- CP-element group 780: 	795 
    -- CP-element group 780:  members (3) 
      -- CP-element group 780: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Sample/ack
      -- CP-element group 780: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Sample/$exit
      -- CP-element group 780: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_sample_complete
      -- 
    ack_11104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 780_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5107_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(780)); -- 
    -- CP-element group 781:  transition  input  output  bypass 
    -- CP-element group 781: predecessors 
    -- CP-element group 781: 	760 
    -- CP-element group 781: successors 
    -- CP-element group 781: 	782 
    -- CP-element group 781:  members (11) 
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_base_plus_offset/sum_rename_ack
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_request/$entry
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_sample_start_
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_request/req
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_root_address_calculated
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_base_plus_offset/sum_rename_req
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_base_plus_offset/$exit
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_base_plus_offset/$entry
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Update/ack
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_final_index_sum_regn_Update/$exit
      -- CP-element group 781: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5107_offset_calculated
      -- 
    ack_11109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 781_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5107_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(781)); -- 
    req_11118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(781), ack => addr_of_5108_final_reg_req_0); -- 
    -- CP-element group 782:  transition  input  bypass 
    -- CP-element group 782: predecessors 
    -- CP-element group 782: 	781 
    -- CP-element group 782: successors 
    -- CP-element group 782:  members (3) 
      -- CP-element group 782: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_request/$exit
      -- CP-element group 782: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_sample_completed_
      -- CP-element group 782: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_request/ack
      -- 
    ack_11119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 782_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5108_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(782)); -- 
    -- CP-element group 783:  join  fork  transition  input  output  bypass 
    -- CP-element group 783: predecessors 
    -- CP-element group 783: 	760 
    -- CP-element group 783: successors 
    -- CP-element group 783: 	784 
    -- CP-element group 783:  members (24) 
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/word_access_start/word_0/$entry
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/word_access_start/word_0/rr
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_update_completed_
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/word_access_start/$entry
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/$entry
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_word_addrgen/root_register_ack
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_word_addrgen/root_register_req
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_word_addrgen/$exit
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_word_addrgen/$entry
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_plus_offset/sum_rename_ack
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_plus_offset/sum_rename_req
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_plus_offset/$exit
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_plus_offset/$entry
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_addr_resize/base_resize_ack
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_addr_resize/base_resize_req
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_addr_resize/$exit
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_addr_resize/$entry
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_address_resized
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_root_address_calculated
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_word_address_calculated
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_base_address_calculated
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_sample_start_
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_complete/ack
      -- CP-element group 783: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5108_complete/$exit
      -- 
    ack_11124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 783_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5108_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(783)); -- 
    rr_11157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(783), ack => ptr_deref_5112_load_0_req_0); -- 
    -- CP-element group 784:  transition  input  bypass 
    -- CP-element group 784: predecessors 
    -- CP-element group 784: 	783 
    -- CP-element group 784: successors 
    -- CP-element group 784:  members (5) 
      -- CP-element group 784: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/word_access_start/$exit
      -- CP-element group 784: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/word_access_start/word_0/$exit
      -- CP-element group 784: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/word_access_start/word_0/ra
      -- CP-element group 784: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Sample/$exit
      -- CP-element group 784: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_sample_completed_
      -- 
    ra_11158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 784_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5112_load_0_ack_0, ack => zeropad3D_CP_2152_elements(784)); -- 
    -- CP-element group 785:  transition  input  bypass 
    -- CP-element group 785: predecessors 
    -- CP-element group 785: 	760 
    -- CP-element group 785: successors 
    -- CP-element group 785: 	792 
    -- CP-element group 785:  members (9) 
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/$exit
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/word_access_complete/$exit
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/word_access_complete/word_0/$exit
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/word_access_complete/word_0/ca
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/ptr_deref_5112_Merge/$entry
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/ptr_deref_5112_Merge/$exit
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/ptr_deref_5112_Merge/merge_req
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_update_completed_
      -- CP-element group 785: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5112_Update/ptr_deref_5112_Merge/merge_ack
      -- 
    ca_11169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 785_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5112_load_0_ack_1, ack => zeropad3D_CP_2152_elements(785)); -- 
    -- CP-element group 786:  transition  input  bypass 
    -- CP-element group 786: predecessors 
    -- CP-element group 786: 	777 
    -- CP-element group 786: successors 
    -- CP-element group 786:  members (3) 
      -- CP-element group 786: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Sample/ra
      -- CP-element group 786: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Sample/$exit
      -- CP-element group 786: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_sample_completed_
      -- 
    ra_11183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 786_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5126_inst_ack_0, ack => zeropad3D_CP_2152_elements(786)); -- 
    -- CP-element group 787:  transition  input  output  bypass 
    -- CP-element group 787: predecessors 
    -- CP-element group 787: 	760 
    -- CP-element group 787: successors 
    -- CP-element group 787: 	788 
    -- CP-element group 787:  members (16) 
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_resize_1/$entry
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_resize_1/$exit
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_resize_1/index_resize_req
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_resize_1/index_resize_ack
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_scale_1/$entry
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_scale_1/$exit
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_scale_1/scale_rename_req
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_scale_1/scale_rename_ack
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_computed_1
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_scaled_1
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_index_resized_1
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Sample/req
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Update/ca
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_Update/$exit
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Sample/$entry
      -- CP-element group 787: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/type_cast_5126_update_completed_
      -- 
    ca_11188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 787_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5126_inst_ack_1, ack => zeropad3D_CP_2152_elements(787)); -- 
    req_11213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(787), ack => array_obj_ref_5132_index_offset_req_0); -- 
    -- CP-element group 788:  transition  input  bypass 
    -- CP-element group 788: predecessors 
    -- CP-element group 788: 	787 
    -- CP-element group 788: successors 
    -- CP-element group 788: 	795 
    -- CP-element group 788:  members (3) 
      -- CP-element group 788: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Sample/ack
      -- CP-element group 788: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Sample/$exit
      -- CP-element group 788: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_sample_complete
      -- 
    ack_11214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 788_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5132_index_offset_ack_0, ack => zeropad3D_CP_2152_elements(788)); -- 
    -- CP-element group 789:  transition  input  output  bypass 
    -- CP-element group 789: predecessors 
    -- CP-element group 789: 	760 
    -- CP-element group 789: successors 
    -- CP-element group 789: 	790 
    -- CP-element group 789:  members (11) 
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Update/$exit
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_base_plus_offset/$entry
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_final_index_sum_regn_Update/ack
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_base_plus_offset/$exit
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_offset_calculated
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_root_address_calculated
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_sample_start_
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_request/$entry
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_request/req
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_base_plus_offset/sum_rename_ack
      -- CP-element group 789: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/array_obj_ref_5132_base_plus_offset/sum_rename_req
      -- 
    ack_11219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 789_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_5132_index_offset_ack_1, ack => zeropad3D_CP_2152_elements(789)); -- 
    req_11228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_11228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(789), ack => addr_of_5133_final_reg_req_0); -- 
    -- CP-element group 790:  transition  input  bypass 
    -- CP-element group 790: predecessors 
    -- CP-element group 790: 	789 
    -- CP-element group 790: successors 
    -- CP-element group 790:  members (3) 
      -- CP-element group 790: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_sample_completed_
      -- CP-element group 790: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_request/ack
      -- CP-element group 790: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_request/$exit
      -- 
    ack_11229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 790_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5133_final_reg_ack_0, ack => zeropad3D_CP_2152_elements(790)); -- 
    -- CP-element group 791:  fork  transition  input  bypass 
    -- CP-element group 791: predecessors 
    -- CP-element group 791: 	760 
    -- CP-element group 791: successors 
    -- CP-element group 791: 	792 
    -- CP-element group 791:  members (19) 
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_word_addrgen/$exit
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_word_addrgen/root_register_req
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_word_addrgen/root_register_ack
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_update_completed_
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_plus_offset/sum_rename_ack
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_plus_offset/sum_rename_req
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_plus_offset/$exit
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_plus_offset/$entry
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_addr_resize/base_resize_ack
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_addr_resize/base_resize_req
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_addr_resize/$exit
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_addr_resize/$entry
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_address_resized
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_root_address_calculated
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_word_address_calculated
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_base_address_calculated
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_complete/ack
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/addr_of_5133_complete/$exit
      -- CP-element group 791: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_word_addrgen/$entry
      -- 
    ack_11234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 791_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_5133_final_reg_ack_1, ack => zeropad3D_CP_2152_elements(791)); -- 
    -- CP-element group 792:  join  transition  output  bypass 
    -- CP-element group 792: predecessors 
    -- CP-element group 792: 	785 
    -- CP-element group 792: 	791 
    -- CP-element group 792: successors 
    -- CP-element group 792: 	793 
    -- CP-element group 792:  members (9) 
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/ptr_deref_5136_Split/$exit
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/ptr_deref_5136_Split/split_req
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/ptr_deref_5136_Split/split_ack
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/word_access_start/word_0/$entry
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/word_access_start/$entry
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/ptr_deref_5136_Split/$entry
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/$entry
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_sample_start_
      -- CP-element group 792: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/word_access_start/word_0/rr
      -- 
    rr_11272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(792), ack => ptr_deref_5136_store_0_req_0); -- 
    zeropad3D_cp_element_group_792: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_792"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(785) & zeropad3D_CP_2152_elements(791);
      gj_zeropad3D_cp_element_group_792 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(792), clk => clk, reset => reset); --
    end block;
    -- CP-element group 793:  transition  input  bypass 
    -- CP-element group 793: predecessors 
    -- CP-element group 793: 	792 
    -- CP-element group 793: successors 
    -- CP-element group 793:  members (5) 
      -- CP-element group 793: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/$exit
      -- CP-element group 793: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_sample_completed_
      -- CP-element group 793: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/word_access_start/word_0/ra
      -- CP-element group 793: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/word_access_start/word_0/$exit
      -- CP-element group 793: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Sample/word_access_start/$exit
      -- 
    ra_11273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 793_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5136_store_0_ack_0, ack => zeropad3D_CP_2152_elements(793)); -- 
    -- CP-element group 794:  transition  input  bypass 
    -- CP-element group 794: predecessors 
    -- CP-element group 794: 	760 
    -- CP-element group 794: successors 
    -- CP-element group 794: 	795 
    -- CP-element group 794:  members (5) 
      -- CP-element group 794: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/word_access_complete/word_0/$exit
      -- CP-element group 794: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/word_access_complete/word_0/ca
      -- CP-element group 794: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/word_access_complete/$exit
      -- CP-element group 794: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_update_completed_
      -- CP-element group 794: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/ptr_deref_5136_Update/$exit
      -- 
    ca_11284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 794_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_5136_store_0_ack_1, ack => zeropad3D_CP_2152_elements(794)); -- 
    -- CP-element group 795:  join  transition  place  bypass 
    -- CP-element group 795: predecessors 
    -- CP-element group 795: 	780 
    -- CP-element group 795: 	788 
    -- CP-element group 795: 	794 
    -- CP-element group 795: successors 
    -- CP-element group 795: 	1168 
    -- CP-element group 795:  members (5) 
      -- CP-element group 795: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138__exit__
      -- CP-element group 795: 	 branch_block_stmt_714/ifx_xelse1617_ifx_xend1665
      -- CP-element group 795: 	 branch_block_stmt_714/assign_stmt_5038_to_assign_stmt_5138/$exit
      -- CP-element group 795: 	 branch_block_stmt_714/ifx_xelse1617_ifx_xend1665_PhiReq/$entry
      -- CP-element group 795: 	 branch_block_stmt_714/ifx_xelse1617_ifx_xend1665_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_795: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_795"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(780) & zeropad3D_CP_2152_elements(788) & zeropad3D_CP_2152_elements(794);
      gj_zeropad3D_cp_element_group_795 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(795), clk => clk, reset => reset); --
    end block;
    -- CP-element group 796:  transition  input  bypass 
    -- CP-element group 796: predecessors 
    -- CP-element group 796: 	1168 
    -- CP-element group 796: successors 
    -- CP-element group 796:  members (3) 
      -- CP-element group 796: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Sample/ra
      -- CP-element group 796: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Sample/$exit
      -- CP-element group 796: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_sample_completed_
      -- 
    ra_11296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 796_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5144_inst_ack_0, ack => zeropad3D_CP_2152_elements(796)); -- 
    -- CP-element group 797:  branch  transition  place  input  output  bypass 
    -- CP-element group 797: predecessors 
    -- CP-element group 797: 	1168 
    -- CP-element group 797: successors 
    -- CP-element group 797: 	798 
    -- CP-element group 797: 	799 
    -- CP-element group 797:  members (13) 
      -- CP-element group 797: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158__exit__
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159__entry__
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159_eval_test/$entry
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159_dead_link/$entry
      -- CP-element group 797: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Update/ca
      -- CP-element group 797: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Update/$exit
      -- CP-element group 797: 	 branch_block_stmt_714/R_cmp1673_5160_place
      -- CP-element group 797: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_update_completed_
      -- CP-element group 797: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/$exit
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159_eval_test/$exit
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159_eval_test/branch_req
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159_if_link/$entry
      -- CP-element group 797: 	 branch_block_stmt_714/if_stmt_5159_else_link/$entry
      -- 
    ca_11301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 797_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5144_inst_ack_1, ack => zeropad3D_CP_2152_elements(797)); -- 
    branch_req_11309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(797), ack => if_stmt_5159_branch_req_0); -- 
    -- CP-element group 798:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 798: predecessors 
    -- CP-element group 798: 	797 
    -- CP-element group 798: successors 
    -- CP-element group 798: 	1177 
    -- CP-element group 798: 	1178 
    -- CP-element group 798: 	1180 
    -- CP-element group 798: 	1181 
    -- CP-element group 798: 	1183 
    -- CP-element group 798: 	1184 
    -- CP-element group 798:  members (40) 
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_5165__exit__
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_5171__entry__
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_5171__exit__
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xend1665_ifx_xthen1675
      -- CP-element group 798: 	 branch_block_stmt_714/if_stmt_5159_if_link/$exit
      -- CP-element group 798: 	 branch_block_stmt_714/if_stmt_5159_if_link/if_choice_transition
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_5171/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/assign_stmt_5171/$exit
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xend1665_ifx_xthen1675_PhiReq/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xend1665_ifx_xthen1675_PhiReq/$exit
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_5165_PhiReqMerge
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_5165_PhiAck/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_5165_PhiAck/$exit
      -- CP-element group 798: 	 branch_block_stmt_714/merge_stmt_5165_PhiAck/dummy
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Sample/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Sample/rr
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Update/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Update/cr
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Sample/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Sample/rr
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Update/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Update/cr
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Sample/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Sample/rr
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Update/$entry
      -- CP-element group 798: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Update/cr
      -- 
    if_choice_transition_11314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 798_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5159_branch_ack_1, ack => zeropad3D_CP_2152_elements(798)); -- 
    rr_14380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_5252_inst_req_0); -- 
    cr_14385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_5252_inst_req_1); -- 
    rr_14403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_5256_inst_req_0); -- 
    cr_14408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_5256_inst_req_1); -- 
    rr_14426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_5262_inst_req_0); -- 
    cr_14431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(798), ack => type_cast_5262_inst_req_1); -- 
    -- CP-element group 799:  fork  transition  place  input  output  bypass 
    -- CP-element group 799: predecessors 
    -- CP-element group 799: 	797 
    -- CP-element group 799: successors 
    -- CP-element group 799: 	800 
    -- CP-element group 799: 	801 
    -- CP-element group 799: 	802 
    -- CP-element group 799: 	803 
    -- CP-element group 799: 	805 
    -- CP-element group 799: 	808 
    -- CP-element group 799: 	810 
    -- CP-element group 799: 	811 
    -- CP-element group 799: 	812 
    -- CP-element group 799: 	814 
    -- CP-element group 799:  members (54) 
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_5173__exit__
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238__entry__
      -- CP-element group 799: 	 branch_block_stmt_714/ifx_xend1665_ifx_xelse1680
      -- CP-element group 799: 	 branch_block_stmt_714/if_stmt_5159_else_link/$exit
      -- CP-element group 799: 	 branch_block_stmt_714/if_stmt_5159_else_link/else_choice_transition
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_sample_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Sample/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Sample/rr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_sample_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_word_address_calculated
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_root_address_calculated
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/word_access_start/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/word_access_start/word_0/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/word_access_start/word_0/rr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/word_access_complete/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/word_access_complete/word_0/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/word_access_complete/word_0/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_sample_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_word_address_calculated
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_root_address_calculated
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/word_access_start/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/word_access_start/word_0/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/word_access_start/word_0/rr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/word_access_complete/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/word_access_complete/word_0/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/word_access_complete/word_0/cr
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_update_start_
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Update/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Update/cr
      -- CP-element group 799: 	 branch_block_stmt_714/ifx_xend1665_ifx_xelse1680_PhiReq/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/ifx_xend1665_ifx_xelse1680_PhiReq/$exit
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_5173_PhiReqMerge
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_5173_PhiAck/$entry
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_5173_PhiAck/$exit
      -- CP-element group 799: 	 branch_block_stmt_714/merge_stmt_5173_PhiAck/dummy
      -- 
    else_choice_transition_11318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 799_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5159_branch_ack_0, ack => zeropad3D_CP_2152_elements(799)); -- 
    rr_11334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_5183_inst_req_0); -- 
    cr_11339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_5183_inst_req_1); -- 
    rr_11356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => LOAD_col_high_5186_load_0_req_0); -- 
    cr_11367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => LOAD_col_high_5186_load_0_req_1); -- 
    cr_11386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_5190_inst_req_1); -- 
    cr_11400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_5204_inst_req_1); -- 
    cr_11414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_5220_inst_req_1); -- 
    rr_11431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => LOAD_row_high_5223_load_0_req_0); -- 
    cr_11442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => LOAD_row_high_5223_load_0_req_1); -- 
    cr_11461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(799), ack => type_cast_5227_inst_req_1); -- 
    -- CP-element group 800:  transition  input  bypass 
    -- CP-element group 800: predecessors 
    -- CP-element group 800: 	799 
    -- CP-element group 800: successors 
    -- CP-element group 800:  members (3) 
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_sample_completed_
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Sample/$exit
      -- CP-element group 800: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Sample/ra
      -- 
    ra_11335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 800_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5183_inst_ack_0, ack => zeropad3D_CP_2152_elements(800)); -- 
    -- CP-element group 801:  transition  input  bypass 
    -- CP-element group 801: predecessors 
    -- CP-element group 801: 	799 
    -- CP-element group 801: successors 
    -- CP-element group 801: 	806 
    -- CP-element group 801:  members (3) 
      -- CP-element group 801: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_update_completed_
      -- CP-element group 801: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Update/$exit
      -- CP-element group 801: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5183_Update/ca
      -- 
    ca_11340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 801_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5183_inst_ack_1, ack => zeropad3D_CP_2152_elements(801)); -- 
    -- CP-element group 802:  transition  input  bypass 
    -- CP-element group 802: predecessors 
    -- CP-element group 802: 	799 
    -- CP-element group 802: successors 
    -- CP-element group 802:  members (5) 
      -- CP-element group 802: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_sample_completed_
      -- CP-element group 802: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/$exit
      -- CP-element group 802: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/word_access_start/$exit
      -- CP-element group 802: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/word_access_start/word_0/$exit
      -- CP-element group 802: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Sample/word_access_start/word_0/ra
      -- 
    ra_11357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 802_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_5186_load_0_ack_0, ack => zeropad3D_CP_2152_elements(802)); -- 
    -- CP-element group 803:  transition  input  output  bypass 
    -- CP-element group 803: predecessors 
    -- CP-element group 803: 	799 
    -- CP-element group 803: successors 
    -- CP-element group 803: 	804 
    -- CP-element group 803:  members (12) 
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_update_completed_
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/word_access_complete/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/word_access_complete/word_0/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/word_access_complete/word_0/ca
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/LOAD_col_high_5186_Merge/$entry
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/LOAD_col_high_5186_Merge/$exit
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/LOAD_col_high_5186_Merge/merge_req
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_col_high_5186_Update/LOAD_col_high_5186_Merge/merge_ack
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_sample_start_
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Sample/$entry
      -- CP-element group 803: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Sample/rr
      -- 
    ca_11368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 803_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_col_high_5186_load_0_ack_1, ack => zeropad3D_CP_2152_elements(803)); -- 
    rr_11381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(803), ack => type_cast_5190_inst_req_0); -- 
    -- CP-element group 804:  transition  input  bypass 
    -- CP-element group 804: predecessors 
    -- CP-element group 804: 	803 
    -- CP-element group 804: successors 
    -- CP-element group 804:  members (3) 
      -- CP-element group 804: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_sample_completed_
      -- CP-element group 804: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Sample/$exit
      -- CP-element group 804: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Sample/ra
      -- 
    ra_11382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 804_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5190_inst_ack_0, ack => zeropad3D_CP_2152_elements(804)); -- 
    -- CP-element group 805:  transition  input  bypass 
    -- CP-element group 805: predecessors 
    -- CP-element group 805: 	799 
    -- CP-element group 805: successors 
    -- CP-element group 805: 	806 
    -- CP-element group 805:  members (3) 
      -- CP-element group 805: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_update_completed_
      -- CP-element group 805: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Update/$exit
      -- CP-element group 805: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5190_Update/ca
      -- 
    ca_11387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 805_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5190_inst_ack_1, ack => zeropad3D_CP_2152_elements(805)); -- 
    -- CP-element group 806:  join  transition  output  bypass 
    -- CP-element group 806: predecessors 
    -- CP-element group 806: 	801 
    -- CP-element group 806: 	805 
    -- CP-element group 806: successors 
    -- CP-element group 806: 	807 
    -- CP-element group 806:  members (3) 
      -- CP-element group 806: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_sample_start_
      -- CP-element group 806: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Sample/$entry
      -- CP-element group 806: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Sample/rr
      -- 
    rr_11395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(806), ack => type_cast_5204_inst_req_0); -- 
    zeropad3D_cp_element_group_806: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_806"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(801) & zeropad3D_CP_2152_elements(805);
      gj_zeropad3D_cp_element_group_806 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(806), clk => clk, reset => reset); --
    end block;
    -- CP-element group 807:  transition  input  bypass 
    -- CP-element group 807: predecessors 
    -- CP-element group 807: 	806 
    -- CP-element group 807: successors 
    -- CP-element group 807:  members (3) 
      -- CP-element group 807: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_sample_completed_
      -- CP-element group 807: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Sample/$exit
      -- CP-element group 807: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Sample/ra
      -- 
    ra_11396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 807_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5204_inst_ack_0, ack => zeropad3D_CP_2152_elements(807)); -- 
    -- CP-element group 808:  transition  input  output  bypass 
    -- CP-element group 808: predecessors 
    -- CP-element group 808: 	799 
    -- CP-element group 808: successors 
    -- CP-element group 808: 	809 
    -- CP-element group 808:  members (6) 
      -- CP-element group 808: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_update_completed_
      -- CP-element group 808: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Update/$exit
      -- CP-element group 808: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5204_Update/ca
      -- CP-element group 808: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_sample_start_
      -- CP-element group 808: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Sample/$entry
      -- CP-element group 808: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Sample/rr
      -- 
    ca_11401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 808_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5204_inst_ack_1, ack => zeropad3D_CP_2152_elements(808)); -- 
    rr_11409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(808), ack => type_cast_5220_inst_req_0); -- 
    -- CP-element group 809:  transition  input  bypass 
    -- CP-element group 809: predecessors 
    -- CP-element group 809: 	808 
    -- CP-element group 809: successors 
    -- CP-element group 809:  members (3) 
      -- CP-element group 809: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_sample_completed_
      -- CP-element group 809: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Sample/$exit
      -- CP-element group 809: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Sample/ra
      -- 
    ra_11410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 809_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5220_inst_ack_0, ack => zeropad3D_CP_2152_elements(809)); -- 
    -- CP-element group 810:  transition  input  bypass 
    -- CP-element group 810: predecessors 
    -- CP-element group 810: 	799 
    -- CP-element group 810: successors 
    -- CP-element group 810: 	815 
    -- CP-element group 810:  members (3) 
      -- CP-element group 810: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_update_completed_
      -- CP-element group 810: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Update/$exit
      -- CP-element group 810: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5220_Update/ca
      -- 
    ca_11415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 810_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5220_inst_ack_1, ack => zeropad3D_CP_2152_elements(810)); -- 
    -- CP-element group 811:  transition  input  bypass 
    -- CP-element group 811: predecessors 
    -- CP-element group 811: 	799 
    -- CP-element group 811: successors 
    -- CP-element group 811:  members (5) 
      -- CP-element group 811: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_sample_completed_
      -- CP-element group 811: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/word_access_start/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/word_access_start/word_0/$exit
      -- CP-element group 811: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Sample/word_access_start/word_0/ra
      -- 
    ra_11432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 811_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_5223_load_0_ack_0, ack => zeropad3D_CP_2152_elements(811)); -- 
    -- CP-element group 812:  transition  input  output  bypass 
    -- CP-element group 812: predecessors 
    -- CP-element group 812: 	799 
    -- CP-element group 812: successors 
    -- CP-element group 812: 	813 
    -- CP-element group 812:  members (12) 
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_update_completed_
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/$exit
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/word_access_complete/$exit
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/word_access_complete/word_0/$exit
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/word_access_complete/word_0/ca
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/LOAD_row_high_5223_Merge/$entry
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/LOAD_row_high_5223_Merge/$exit
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/LOAD_row_high_5223_Merge/merge_req
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/LOAD_row_high_5223_Update/LOAD_row_high_5223_Merge/merge_ack
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_sample_start_
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Sample/$entry
      -- CP-element group 812: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Sample/rr
      -- 
    ca_11443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 812_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_row_high_5223_load_0_ack_1, ack => zeropad3D_CP_2152_elements(812)); -- 
    rr_11456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(812), ack => type_cast_5227_inst_req_0); -- 
    -- CP-element group 813:  transition  input  bypass 
    -- CP-element group 813: predecessors 
    -- CP-element group 813: 	812 
    -- CP-element group 813: successors 
    -- CP-element group 813:  members (3) 
      -- CP-element group 813: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_sample_completed_
      -- CP-element group 813: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Sample/$exit
      -- CP-element group 813: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Sample/ra
      -- 
    ra_11457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 813_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5227_inst_ack_0, ack => zeropad3D_CP_2152_elements(813)); -- 
    -- CP-element group 814:  transition  input  bypass 
    -- CP-element group 814: predecessors 
    -- CP-element group 814: 	799 
    -- CP-element group 814: successors 
    -- CP-element group 814: 	815 
    -- CP-element group 814:  members (3) 
      -- CP-element group 814: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_update_completed_
      -- CP-element group 814: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Update/$exit
      -- CP-element group 814: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/type_cast_5227_Update/ca
      -- 
    ca_11462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 814_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5227_inst_ack_1, ack => zeropad3D_CP_2152_elements(814)); -- 
    -- CP-element group 815:  branch  join  transition  place  output  bypass 
    -- CP-element group 815: predecessors 
    -- CP-element group 815: 	810 
    -- CP-element group 815: 	814 
    -- CP-element group 815: successors 
    -- CP-element group 815: 	816 
    -- CP-element group 815: 	817 
    -- CP-element group 815:  members (10) 
      -- CP-element group 815: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238__exit__
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239__entry__
      -- CP-element group 815: 	 branch_block_stmt_714/assign_stmt_5179_to_assign_stmt_5238/$exit
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239_dead_link/$entry
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239_eval_test/$entry
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239_eval_test/$exit
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239_eval_test/branch_req
      -- CP-element group 815: 	 branch_block_stmt_714/R_cmp1706_5240_place
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239_if_link/$entry
      -- CP-element group 815: 	 branch_block_stmt_714/if_stmt_5239_else_link/$entry
      -- 
    branch_req_11470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_11470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(815), ack => if_stmt_5239_branch_req_0); -- 
    zeropad3D_cp_element_group_815: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_815"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(810) & zeropad3D_CP_2152_elements(814);
      gj_zeropad3D_cp_element_group_815 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(815), clk => clk, reset => reset); --
    end block;
    -- CP-element group 816:  fork  transition  place  input  output  bypass 
    -- CP-element group 816: predecessors 
    -- CP-element group 816: 	815 
    -- CP-element group 816: successors 
    -- CP-element group 816: 	818 
    -- CP-element group 816: 	819 
    -- CP-element group 816:  members (18) 
      -- CP-element group 816: 	 branch_block_stmt_714/merge_stmt_5267__exit__
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270__entry__
      -- CP-element group 816: 	 branch_block_stmt_714/if_stmt_5239_if_link/$exit
      -- CP-element group 816: 	 branch_block_stmt_714/if_stmt_5239_if_link/if_choice_transition
      -- CP-element group 816: 	 branch_block_stmt_714/ifx_xelse1680_whilex_xend1716
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/$entry
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_sample_start_
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_update_start_
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/$entry
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/crr
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/$entry
      -- CP-element group 816: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/ccr
      -- CP-element group 816: 	 branch_block_stmt_714/ifx_xelse1680_whilex_xend1716_PhiReq/$entry
      -- CP-element group 816: 	 branch_block_stmt_714/ifx_xelse1680_whilex_xend1716_PhiReq/$exit
      -- CP-element group 816: 	 branch_block_stmt_714/merge_stmt_5267_PhiReqMerge
      -- CP-element group 816: 	 branch_block_stmt_714/merge_stmt_5267_PhiAck/$entry
      -- CP-element group 816: 	 branch_block_stmt_714/merge_stmt_5267_PhiAck/$exit
      -- CP-element group 816: 	 branch_block_stmt_714/merge_stmt_5267_PhiAck/dummy
      -- 
    if_choice_transition_11475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 816_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5239_branch_ack_1, ack => zeropad3D_CP_2152_elements(816)); -- 
    crr_11492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_11492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(816), ack => call_stmt_5270_call_req_0); -- 
    ccr_11497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_11497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(816), ack => call_stmt_5270_call_req_1); -- 
    -- CP-element group 817:  fork  transition  place  input  output  bypass 
    -- CP-element group 817: predecessors 
    -- CP-element group 817: 	815 
    -- CP-element group 817: successors 
    -- CP-element group 817: 	1169 
    -- CP-element group 817: 	1170 
    -- CP-element group 817: 	1171 
    -- CP-element group 817: 	1173 
    -- CP-element group 817: 	1174 
    -- CP-element group 817:  members (22) 
      -- CP-element group 817: 	 branch_block_stmt_714/if_stmt_5239_else_link/$exit
      -- CP-element group 817: 	 branch_block_stmt_714/if_stmt_5239_else_link/else_choice_transition
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5246/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Sample/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Sample/rr
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Update/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Update/cr
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Sample/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Sample/rr
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Update/$entry
      -- CP-element group 817: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Update/cr
      -- 
    else_choice_transition_11479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 817_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_5239_branch_ack_0, ack => zeropad3D_CP_2152_elements(817)); -- 
    rr_14331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(817), ack => type_cast_5258_inst_req_0); -- 
    cr_14336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(817), ack => type_cast_5258_inst_req_1); -- 
    rr_14354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_14354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(817), ack => type_cast_5264_inst_req_0); -- 
    cr_14359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_14359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(817), ack => type_cast_5264_inst_req_1); -- 
    -- CP-element group 818:  transition  input  bypass 
    -- CP-element group 818: predecessors 
    -- CP-element group 818: 	816 
    -- CP-element group 818: successors 
    -- CP-element group 818:  members (3) 
      -- CP-element group 818: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_sample_completed_
      -- CP-element group 818: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/$exit
      -- CP-element group 818: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Sample/cra
      -- 
    cra_11493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 818_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_5270_call_ack_0, ack => zeropad3D_CP_2152_elements(818)); -- 
    -- CP-element group 819:  transition  place  input  bypass 
    -- CP-element group 819: predecessors 
    -- CP-element group 819: 	816 
    -- CP-element group 819: successors 
    -- CP-element group 819:  members (16) 
      -- CP-element group 819: 	 branch_block_stmt_714/branch_block_stmt_714__exit__
      -- CP-element group 819: 	 branch_block_stmt_714/$exit
      -- CP-element group 819: 	 $exit
      -- CP-element group 819: 	 branch_block_stmt_714/call_stmt_5270__exit__
      -- CP-element group 819: 	 branch_block_stmt_714/return__
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_5272__exit__
      -- CP-element group 819: 	 branch_block_stmt_714/call_stmt_5270/$exit
      -- CP-element group 819: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_update_completed_
      -- CP-element group 819: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/$exit
      -- CP-element group 819: 	 branch_block_stmt_714/call_stmt_5270/call_stmt_5270_Update/cca
      -- CP-element group 819: 	 branch_block_stmt_714/return___PhiReq/$entry
      -- CP-element group 819: 	 branch_block_stmt_714/return___PhiReq/$exit
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_5272_PhiReqMerge
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_5272_PhiAck/$entry
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_5272_PhiAck/$exit
      -- CP-element group 819: 	 branch_block_stmt_714/merge_stmt_5272_PhiAck/dummy
      -- 
    cca_11498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 819_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_5270_call_ack_1, ack => zeropad3D_CP_2152_elements(819)); -- 
    -- CP-element group 820:  transition  output  delay-element  bypass 
    -- CP-element group 820: predecessors 
    -- CP-element group 820: 	58 
    -- CP-element group 820: successors 
    -- CP-element group 820: 	823 
    -- CP-element group 820:  members (4) 
      -- CP-element group 820: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/$exit
      -- CP-element group 820: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$exit
      -- CP-element group 820: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_903_konst_delay_trans
      -- CP-element group 820: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_req
      -- 
    phi_stmt_899_req_11509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_899_req_11509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(820), ack => phi_stmt_899_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(820) is a control-delay.
    cp_element_820_delay: control_delay_element  generic map(name => " 820_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(58), ack => zeropad3D_CP_2152_elements(820), clk => clk, reset =>reset);
    -- CP-element group 821:  transition  output  delay-element  bypass 
    -- CP-element group 821: predecessors 
    -- CP-element group 821: 	58 
    -- CP-element group 821: successors 
    -- CP-element group 821: 	823 
    -- CP-element group 821:  members (4) 
      -- CP-element group 821: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/$exit
      -- CP-element group 821: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$exit
      -- CP-element group 821: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_910_konst_delay_trans
      -- CP-element group 821: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_req
      -- 
    phi_stmt_906_req_11517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_906_req_11517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(821), ack => phi_stmt_906_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(821) is a control-delay.
    cp_element_821_delay: control_delay_element  generic map(name => " 821_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(58), ack => zeropad3D_CP_2152_elements(821), clk => clk, reset =>reset);
    -- CP-element group 822:  transition  output  delay-element  bypass 
    -- CP-element group 822: predecessors 
    -- CP-element group 822: 	58 
    -- CP-element group 822: successors 
    -- CP-element group 822: 	823 
    -- CP-element group 822:  members (4) 
      -- CP-element group 822: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/$exit
      -- CP-element group 822: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$exit
      -- CP-element group 822: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_917_konst_delay_trans
      -- CP-element group 822: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_req
      -- 
    phi_stmt_913_req_11525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_913_req_11525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(822), ack => phi_stmt_913_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(822) is a control-delay.
    cp_element_822_delay: control_delay_element  generic map(name => " 822_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(58), ack => zeropad3D_CP_2152_elements(822), clk => clk, reset =>reset);
    -- CP-element group 823:  join  transition  bypass 
    -- CP-element group 823: predecessors 
    -- CP-element group 823: 	820 
    -- CP-element group 823: 	821 
    -- CP-element group 823: 	822 
    -- CP-element group 823: successors 
    -- CP-element group 823: 	834 
    -- CP-element group 823:  members (1) 
      -- CP-element group 823: 	 branch_block_stmt_714/entry_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_823: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_823"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(820) & zeropad3D_CP_2152_elements(821) & zeropad3D_CP_2152_elements(822);
      gj_zeropad3D_cp_element_group_823 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(823), clk => clk, reset => reset); --
    end block;
    -- CP-element group 824:  transition  input  bypass 
    -- CP-element group 824: predecessors 
    -- CP-element group 824: 	1 
    -- CP-element group 824: successors 
    -- CP-element group 824: 	826 
    -- CP-element group 824:  members (2) 
      -- CP-element group 824: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/$exit
      -- CP-element group 824: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Sample/ra
      -- 
    ra_11545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 824_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => zeropad3D_CP_2152_elements(824)); -- 
    -- CP-element group 825:  transition  input  bypass 
    -- CP-element group 825: predecessors 
    -- CP-element group 825: 	1 
    -- CP-element group 825: successors 
    -- CP-element group 825: 	826 
    -- CP-element group 825:  members (2) 
      -- CP-element group 825: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/$exit
      -- CP-element group 825: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/Update/ca
      -- 
    ca_11550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 825_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => zeropad3D_CP_2152_elements(825)); -- 
    -- CP-element group 826:  join  transition  output  bypass 
    -- CP-element group 826: predecessors 
    -- CP-element group 826: 	824 
    -- CP-element group 826: 	825 
    -- CP-element group 826: successors 
    -- CP-element group 826: 	833 
    -- CP-element group 826:  members (5) 
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_sources/type_cast_905/SplitProtocol/$exit
      -- CP-element group 826: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_899/phi_stmt_899_req
      -- 
    phi_stmt_899_req_11551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_899_req_11551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(826), ack => phi_stmt_899_req_1); -- 
    zeropad3D_cp_element_group_826: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_826"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(824) & zeropad3D_CP_2152_elements(825);
      gj_zeropad3D_cp_element_group_826 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(826), clk => clk, reset => reset); --
    end block;
    -- CP-element group 827:  transition  input  bypass 
    -- CP-element group 827: predecessors 
    -- CP-element group 827: 	1 
    -- CP-element group 827: successors 
    -- CP-element group 827: 	829 
    -- CP-element group 827:  members (2) 
      -- CP-element group 827: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/$exit
      -- CP-element group 827: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Sample/ra
      -- 
    ra_11568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 827_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_912_inst_ack_0, ack => zeropad3D_CP_2152_elements(827)); -- 
    -- CP-element group 828:  transition  input  bypass 
    -- CP-element group 828: predecessors 
    -- CP-element group 828: 	1 
    -- CP-element group 828: successors 
    -- CP-element group 828: 	829 
    -- CP-element group 828:  members (2) 
      -- CP-element group 828: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/$exit
      -- CP-element group 828: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/Update/ca
      -- 
    ca_11573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 828_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_912_inst_ack_1, ack => zeropad3D_CP_2152_elements(828)); -- 
    -- CP-element group 829:  join  transition  output  bypass 
    -- CP-element group 829: predecessors 
    -- CP-element group 829: 	827 
    -- CP-element group 829: 	828 
    -- CP-element group 829: successors 
    -- CP-element group 829: 	833 
    -- CP-element group 829:  members (5) 
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_sources/type_cast_912/SplitProtocol/$exit
      -- CP-element group 829: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_906/phi_stmt_906_req
      -- 
    phi_stmt_906_req_11574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_906_req_11574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(829), ack => phi_stmt_906_req_1); -- 
    zeropad3D_cp_element_group_829: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_829"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(827) & zeropad3D_CP_2152_elements(828);
      gj_zeropad3D_cp_element_group_829 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(829), clk => clk, reset => reset); --
    end block;
    -- CP-element group 830:  transition  input  bypass 
    -- CP-element group 830: predecessors 
    -- CP-element group 830: 	1 
    -- CP-element group 830: successors 
    -- CP-element group 830: 	832 
    -- CP-element group 830:  members (2) 
      -- CP-element group 830: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/$exit
      -- CP-element group 830: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Sample/ra
      -- 
    ra_11591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 830_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_919_inst_ack_0, ack => zeropad3D_CP_2152_elements(830)); -- 
    -- CP-element group 831:  transition  input  bypass 
    -- CP-element group 831: predecessors 
    -- CP-element group 831: 	1 
    -- CP-element group 831: successors 
    -- CP-element group 831: 	832 
    -- CP-element group 831:  members (2) 
      -- CP-element group 831: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/$exit
      -- CP-element group 831: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/Update/ca
      -- 
    ca_11596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 831_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_919_inst_ack_1, ack => zeropad3D_CP_2152_elements(831)); -- 
    -- CP-element group 832:  join  transition  output  bypass 
    -- CP-element group 832: predecessors 
    -- CP-element group 832: 	830 
    -- CP-element group 832: 	831 
    -- CP-element group 832: successors 
    -- CP-element group 832: 	833 
    -- CP-element group 832:  members (5) 
      -- CP-element group 832: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/$exit
      -- CP-element group 832: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/$exit
      -- CP-element group 832: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/$exit
      -- CP-element group 832: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_sources/type_cast_919/SplitProtocol/$exit
      -- CP-element group 832: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/phi_stmt_913/phi_stmt_913_req
      -- 
    phi_stmt_913_req_11597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_913_req_11597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(832), ack => phi_stmt_913_req_1); -- 
    zeropad3D_cp_element_group_832: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_832"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(830) & zeropad3D_CP_2152_elements(831);
      gj_zeropad3D_cp_element_group_832 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(832), clk => clk, reset => reset); --
    end block;
    -- CP-element group 833:  join  transition  bypass 
    -- CP-element group 833: predecessors 
    -- CP-element group 833: 	826 
    -- CP-element group 833: 	829 
    -- CP-element group 833: 	832 
    -- CP-element group 833: successors 
    -- CP-element group 833: 	834 
    -- CP-element group 833:  members (1) 
      -- CP-element group 833: 	 branch_block_stmt_714/ifx_xend184_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_833: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_833"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(826) & zeropad3D_CP_2152_elements(829) & zeropad3D_CP_2152_elements(832);
      gj_zeropad3D_cp_element_group_833 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(833), clk => clk, reset => reset); --
    end block;
    -- CP-element group 834:  merge  fork  transition  place  bypass 
    -- CP-element group 834: predecessors 
    -- CP-element group 834: 	823 
    -- CP-element group 834: 	833 
    -- CP-element group 834: successors 
    -- CP-element group 834: 	835 
    -- CP-element group 834: 	836 
    -- CP-element group 834: 	837 
    -- CP-element group 834:  members (2) 
      -- CP-element group 834: 	 branch_block_stmt_714/merge_stmt_898_PhiReqMerge
      -- CP-element group 834: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(834) <= OrReduce(zeropad3D_CP_2152_elements(823) & zeropad3D_CP_2152_elements(833));
    -- CP-element group 835:  transition  input  bypass 
    -- CP-element group 835: predecessors 
    -- CP-element group 835: 	834 
    -- CP-element group 835: successors 
    -- CP-element group 835: 	838 
    -- CP-element group 835:  members (1) 
      -- CP-element group 835: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/phi_stmt_899_ack
      -- 
    phi_stmt_899_ack_11602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 835_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_899_ack_0, ack => zeropad3D_CP_2152_elements(835)); -- 
    -- CP-element group 836:  transition  input  bypass 
    -- CP-element group 836: predecessors 
    -- CP-element group 836: 	834 
    -- CP-element group 836: successors 
    -- CP-element group 836: 	838 
    -- CP-element group 836:  members (1) 
      -- CP-element group 836: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/phi_stmt_906_ack
      -- 
    phi_stmt_906_ack_11603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 836_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_906_ack_0, ack => zeropad3D_CP_2152_elements(836)); -- 
    -- CP-element group 837:  transition  input  bypass 
    -- CP-element group 837: predecessors 
    -- CP-element group 837: 	834 
    -- CP-element group 837: successors 
    -- CP-element group 837: 	838 
    -- CP-element group 837:  members (1) 
      -- CP-element group 837: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/phi_stmt_913_ack
      -- 
    phi_stmt_913_ack_11604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 837_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_913_ack_0, ack => zeropad3D_CP_2152_elements(837)); -- 
    -- CP-element group 838:  join  fork  transition  place  output  bypass 
    -- CP-element group 838: predecessors 
    -- CP-element group 838: 	835 
    -- CP-element group 838: 	836 
    -- CP-element group 838: 	837 
    -- CP-element group 838: successors 
    -- CP-element group 838: 	59 
    -- CP-element group 838: 	60 
    -- CP-element group 838:  members (10) 
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932__entry__
      -- CP-element group 838: 	 branch_block_stmt_714/merge_stmt_898__exit__
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/$entry
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_sample_start_
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_update_start_
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/$entry
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Sample/rr
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/$entry
      -- CP-element group 838: 	 branch_block_stmt_714/assign_stmt_925_to_assign_stmt_932/type_cast_924_Update/cr
      -- CP-element group 838: 	 branch_block_stmt_714/merge_stmt_898_PhiAck/$exit
      -- 
    rr_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(838), ack => type_cast_924_inst_req_0); -- 
    cr_3171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(838), ack => type_cast_924_inst_req_1); -- 
    zeropad3D_cp_element_group_838: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_838"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(835) & zeropad3D_CP_2152_elements(836) & zeropad3D_CP_2152_elements(837);
      gj_zeropad3D_cp_element_group_838 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(838), clk => clk, reset => reset); --
    end block;
    -- CP-element group 839:  merge  fork  transition  place  output  bypass 
    -- CP-element group 839: predecessors 
    -- CP-element group 839: 	61 
    -- CP-element group 839: 	68 
    -- CP-element group 839: 	71 
    -- CP-element group 839: 	78 
    -- CP-element group 839: successors 
    -- CP-element group 839: 	79 
    -- CP-element group 839: 	80 
    -- CP-element group 839: 	81 
    -- CP-element group 839: 	82 
    -- CP-element group 839: 	85 
    -- CP-element group 839: 	87 
    -- CP-element group 839: 	89 
    -- CP-element group 839: 	91 
    -- CP-element group 839:  members (33) 
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079__entry__
      -- CP-element group 839: 	 branch_block_stmt_714/merge_stmt_1022__exit__
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/cr
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/rr
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_update_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/word_access_complete/word_0/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_update_start
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_sample_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Sample/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_update_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_update_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_Update/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_sample_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/ptr_deref_1076_update_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/cr
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/req
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_Update/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/cr
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/addr_of_1073_complete/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Update/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/req
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/array_obj_ref_1072_final_index_sum_regn_Update/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1026_Sample/rr
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1066_update_start_
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/cr
      -- CP-element group 839: 	 branch_block_stmt_714/assign_stmt_1027_to_assign_stmt_1079/type_cast_1031_Update/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/merge_stmt_1022_PhiReqMerge
      -- CP-element group 839: 	 branch_block_stmt_714/merge_stmt_1022_PhiAck/$entry
      -- CP-element group 839: 	 branch_block_stmt_714/merge_stmt_1022_PhiAck/$exit
      -- CP-element group 839: 	 branch_block_stmt_714/merge_stmt_1022_PhiAck/dummy
      -- 
    cr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => ptr_deref_1076_store_0_req_1); -- 
    rr_3390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => type_cast_1031_inst_req_0); -- 
    cr_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => type_cast_1066_inst_req_1); -- 
    req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => addr_of_1073_final_reg_req_1); -- 
    cr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => type_cast_1026_inst_req_1); -- 
    req_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => array_obj_ref_1072_index_offset_req_1); -- 
    rr_3376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => type_cast_1026_inst_req_0); -- 
    cr_3395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(839), ack => type_cast_1031_inst_req_1); -- 
    zeropad3D_CP_2152_elements(839) <= OrReduce(zeropad3D_CP_2152_elements(61) & zeropad3D_CP_2152_elements(68) & zeropad3D_CP_2152_elements(71) & zeropad3D_CP_2152_elements(78));
    -- CP-element group 840:  merge  fork  transition  place  output  bypass 
    -- CP-element group 840: predecessors 
    -- CP-element group 840: 	92 
    -- CP-element group 840: 	112 
    -- CP-element group 840: successors 
    -- CP-element group 840: 	113 
    -- CP-element group 840: 	114 
    -- CP-element group 840:  members (13) 
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206__entry__
      -- CP-element group 840: 	 branch_block_stmt_714/merge_stmt_1188__exit__
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/$entry
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_sample_start_
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_update_start_
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/$entry
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Sample/rr
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/$entry
      -- CP-element group 840: 	 branch_block_stmt_714/assign_stmt_1193_to_assign_stmt_1206/type_cast_1192_Update/cr
      -- CP-element group 840: 	 branch_block_stmt_714/merge_stmt_1188_PhiReqMerge
      -- CP-element group 840: 	 branch_block_stmt_714/merge_stmt_1188_PhiAck/$entry
      -- CP-element group 840: 	 branch_block_stmt_714/merge_stmt_1188_PhiAck/$exit
      -- CP-element group 840: 	 branch_block_stmt_714/merge_stmt_1188_PhiAck/dummy
      -- 
    rr_3754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(840), ack => type_cast_1192_inst_req_0); -- 
    cr_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(840), ack => type_cast_1192_inst_req_1); -- 
    zeropad3D_CP_2152_elements(840) <= OrReduce(zeropad3D_CP_2152_elements(92) & zeropad3D_CP_2152_elements(112));
    -- CP-element group 841:  transition  input  bypass 
    -- CP-element group 841: predecessors 
    -- CP-element group 841: 	134 
    -- CP-element group 841: successors 
    -- CP-element group 841: 	843 
    -- CP-element group 841:  members (2) 
      -- CP-element group 841: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/$exit
      -- CP-element group 841: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Sample/ra
      -- 
    ra_11724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 841_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_0, ack => zeropad3D_CP_2152_elements(841)); -- 
    -- CP-element group 842:  transition  input  bypass 
    -- CP-element group 842: predecessors 
    -- CP-element group 842: 	134 
    -- CP-element group 842: successors 
    -- CP-element group 842: 	843 
    -- CP-element group 842:  members (2) 
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/$exit
      -- CP-element group 842: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/Update/ca
      -- 
    ca_11729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 842_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_1, ack => zeropad3D_CP_2152_elements(842)); -- 
    -- CP-element group 843:  join  transition  output  bypass 
    -- CP-element group 843: predecessors 
    -- CP-element group 843: 	841 
    -- CP-element group 843: 	842 
    -- CP-element group 843: successors 
    -- CP-element group 843: 	848 
    -- CP-element group 843:  members (5) 
      -- CP-element group 843: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/$exit
      -- CP-element group 843: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$exit
      -- CP-element group 843: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/$exit
      -- CP-element group 843: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1318/SplitProtocol/$exit
      -- CP-element group 843: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_req
      -- 
    phi_stmt_1313_req_11730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1313_req_11730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(843), ack => phi_stmt_1313_req_1); -- 
    zeropad3D_cp_element_group_843: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_843"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(841) & zeropad3D_CP_2152_elements(842);
      gj_zeropad3D_cp_element_group_843 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(843), clk => clk, reset => reset); --
    end block;
    -- CP-element group 844:  transition  output  delay-element  bypass 
    -- CP-element group 844: predecessors 
    -- CP-element group 844: 	134 
    -- CP-element group 844: successors 
    -- CP-element group 844: 	848 
    -- CP-element group 844:  members (4) 
      -- CP-element group 844: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/$exit
      -- CP-element group 844: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$exit
      -- CP-element group 844: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1323_konst_delay_trans
      -- CP-element group 844: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_req
      -- 
    phi_stmt_1319_req_11738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1319_req_11738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(844), ack => phi_stmt_1319_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(844) is a control-delay.
    cp_element_844_delay: control_delay_element  generic map(name => " 844_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(134), ack => zeropad3D_CP_2152_elements(844), clk => clk, reset =>reset);
    -- CP-element group 845:  transition  input  bypass 
    -- CP-element group 845: predecessors 
    -- CP-element group 845: 	134 
    -- CP-element group 845: successors 
    -- CP-element group 845: 	847 
    -- CP-element group 845:  members (2) 
      -- CP-element group 845: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/$exit
      -- CP-element group 845: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Sample/ra
      -- 
    ra_11755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 845_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_0, ack => zeropad3D_CP_2152_elements(845)); -- 
    -- CP-element group 846:  transition  input  bypass 
    -- CP-element group 846: predecessors 
    -- CP-element group 846: 	134 
    -- CP-element group 846: successors 
    -- CP-element group 846: 	847 
    -- CP-element group 846:  members (2) 
      -- CP-element group 846: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/$exit
      -- CP-element group 846: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/Update/ca
      -- 
    ca_11760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 846_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_1, ack => zeropad3D_CP_2152_elements(846)); -- 
    -- CP-element group 847:  join  transition  output  bypass 
    -- CP-element group 847: predecessors 
    -- CP-element group 847: 	845 
    -- CP-element group 847: 	846 
    -- CP-element group 847: successors 
    -- CP-element group 847: 	848 
    -- CP-element group 847:  members (5) 
      -- CP-element group 847: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/$exit
      -- CP-element group 847: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$exit
      -- CP-element group 847: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/$exit
      -- CP-element group 847: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1310/SplitProtocol/$exit
      -- CP-element group 847: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_req
      -- 
    phi_stmt_1307_req_11761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1307_req_11761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(847), ack => phi_stmt_1307_req_0); -- 
    zeropad3D_cp_element_group_847: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_847"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(845) & zeropad3D_CP_2152_elements(846);
      gj_zeropad3D_cp_element_group_847 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(847), clk => clk, reset => reset); --
    end block;
    -- CP-element group 848:  join  transition  bypass 
    -- CP-element group 848: predecessors 
    -- CP-element group 848: 	843 
    -- CP-element group 848: 	844 
    -- CP-element group 848: 	847 
    -- CP-element group 848: successors 
    -- CP-element group 848: 	859 
    -- CP-element group 848:  members (1) 
      -- CP-element group 848: 	 branch_block_stmt_714/ifx_xelse150_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_848: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_848"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(843) & zeropad3D_CP_2152_elements(844) & zeropad3D_CP_2152_elements(847);
      gj_zeropad3D_cp_element_group_848 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(848), clk => clk, reset => reset); --
    end block;
    -- CP-element group 849:  transition  input  bypass 
    -- CP-element group 849: predecessors 
    -- CP-element group 849: 	115 
    -- CP-element group 849: successors 
    -- CP-element group 849: 	851 
    -- CP-element group 849:  members (2) 
      -- CP-element group 849: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/$exit
      -- CP-element group 849: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Sample/ra
      -- 
    ra_11781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 849_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_0, ack => zeropad3D_CP_2152_elements(849)); -- 
    -- CP-element group 850:  transition  input  bypass 
    -- CP-element group 850: predecessors 
    -- CP-element group 850: 	115 
    -- CP-element group 850: successors 
    -- CP-element group 850: 	851 
    -- CP-element group 850:  members (2) 
      -- CP-element group 850: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/$exit
      -- CP-element group 850: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/Update/ca
      -- 
    ca_11786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 850_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_1, ack => zeropad3D_CP_2152_elements(850)); -- 
    -- CP-element group 851:  join  transition  output  bypass 
    -- CP-element group 851: predecessors 
    -- CP-element group 851: 	849 
    -- CP-element group 851: 	850 
    -- CP-element group 851: successors 
    -- CP-element group 851: 	858 
    -- CP-element group 851:  members (5) 
      -- CP-element group 851: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/$exit
      -- CP-element group 851: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/$exit
      -- CP-element group 851: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/$exit
      -- CP-element group 851: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_sources/type_cast_1316/SplitProtocol/$exit
      -- CP-element group 851: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1313/phi_stmt_1313_req
      -- 
    phi_stmt_1313_req_11787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1313_req_11787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(851), ack => phi_stmt_1313_req_0); -- 
    zeropad3D_cp_element_group_851: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_851"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(849) & zeropad3D_CP_2152_elements(850);
      gj_zeropad3D_cp_element_group_851 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(851), clk => clk, reset => reset); --
    end block;
    -- CP-element group 852:  transition  input  bypass 
    -- CP-element group 852: predecessors 
    -- CP-element group 852: 	115 
    -- CP-element group 852: successors 
    -- CP-element group 852: 	854 
    -- CP-element group 852:  members (2) 
      -- CP-element group 852: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/$exit
      -- CP-element group 852: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Sample/ra
      -- 
    ra_11804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 852_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_0, ack => zeropad3D_CP_2152_elements(852)); -- 
    -- CP-element group 853:  transition  input  bypass 
    -- CP-element group 853: predecessors 
    -- CP-element group 853: 	115 
    -- CP-element group 853: successors 
    -- CP-element group 853: 	854 
    -- CP-element group 853:  members (2) 
      -- CP-element group 853: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/$exit
      -- CP-element group 853: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/Update/ca
      -- 
    ca_11809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 853_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_1, ack => zeropad3D_CP_2152_elements(853)); -- 
    -- CP-element group 854:  join  transition  output  bypass 
    -- CP-element group 854: predecessors 
    -- CP-element group 854: 	852 
    -- CP-element group 854: 	853 
    -- CP-element group 854: successors 
    -- CP-element group 854: 	858 
    -- CP-element group 854:  members (5) 
      -- CP-element group 854: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/$exit
      -- CP-element group 854: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/$exit
      -- CP-element group 854: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/$exit
      -- CP-element group 854: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_sources/type_cast_1325/SplitProtocol/$exit
      -- CP-element group 854: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1319/phi_stmt_1319_req
      -- 
    phi_stmt_1319_req_11810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1319_req_11810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(854), ack => phi_stmt_1319_req_1); -- 
    zeropad3D_cp_element_group_854: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_854"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(852) & zeropad3D_CP_2152_elements(853);
      gj_zeropad3D_cp_element_group_854 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(854), clk => clk, reset => reset); --
    end block;
    -- CP-element group 855:  transition  input  bypass 
    -- CP-element group 855: predecessors 
    -- CP-element group 855: 	115 
    -- CP-element group 855: successors 
    -- CP-element group 855: 	857 
    -- CP-element group 855:  members (2) 
      -- CP-element group 855: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/$exit
      -- CP-element group 855: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Sample/ra
      -- 
    ra_11827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 855_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_0, ack => zeropad3D_CP_2152_elements(855)); -- 
    -- CP-element group 856:  transition  input  bypass 
    -- CP-element group 856: predecessors 
    -- CP-element group 856: 	115 
    -- CP-element group 856: successors 
    -- CP-element group 856: 	857 
    -- CP-element group 856:  members (2) 
      -- CP-element group 856: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/$exit
      -- CP-element group 856: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/Update/ca
      -- 
    ca_11832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 856_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_1, ack => zeropad3D_CP_2152_elements(856)); -- 
    -- CP-element group 857:  join  transition  output  bypass 
    -- CP-element group 857: predecessors 
    -- CP-element group 857: 	855 
    -- CP-element group 857: 	856 
    -- CP-element group 857: successors 
    -- CP-element group 857: 	858 
    -- CP-element group 857:  members (5) 
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/$exit
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/$exit
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/$exit
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_sources/type_cast_1312/SplitProtocol/$exit
      -- CP-element group 857: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/phi_stmt_1307/phi_stmt_1307_req
      -- 
    phi_stmt_1307_req_11833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1307_req_11833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(857), ack => phi_stmt_1307_req_1); -- 
    zeropad3D_cp_element_group_857: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_857"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(855) & zeropad3D_CP_2152_elements(856);
      gj_zeropad3D_cp_element_group_857 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(857), clk => clk, reset => reset); --
    end block;
    -- CP-element group 858:  join  transition  bypass 
    -- CP-element group 858: predecessors 
    -- CP-element group 858: 	851 
    -- CP-element group 858: 	854 
    -- CP-element group 858: 	857 
    -- CP-element group 858: successors 
    -- CP-element group 858: 	859 
    -- CP-element group 858:  members (1) 
      -- CP-element group 858: 	 branch_block_stmt_714/ifx_xthen145_ifx_xend184_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_858: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_858"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(851) & zeropad3D_CP_2152_elements(854) & zeropad3D_CP_2152_elements(857);
      gj_zeropad3D_cp_element_group_858 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(858), clk => clk, reset => reset); --
    end block;
    -- CP-element group 859:  merge  fork  transition  place  bypass 
    -- CP-element group 859: predecessors 
    -- CP-element group 859: 	848 
    -- CP-element group 859: 	858 
    -- CP-element group 859: successors 
    -- CP-element group 859: 	860 
    -- CP-element group 859: 	861 
    -- CP-element group 859: 	862 
    -- CP-element group 859:  members (2) 
      -- CP-element group 859: 	 branch_block_stmt_714/merge_stmt_1306_PhiReqMerge
      -- CP-element group 859: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(859) <= OrReduce(zeropad3D_CP_2152_elements(848) & zeropad3D_CP_2152_elements(858));
    -- CP-element group 860:  transition  input  bypass 
    -- CP-element group 860: predecessors 
    -- CP-element group 860: 	859 
    -- CP-element group 860: successors 
    -- CP-element group 860: 	863 
    -- CP-element group 860:  members (1) 
      -- CP-element group 860: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/phi_stmt_1307_ack
      -- 
    phi_stmt_1307_ack_11838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 860_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1307_ack_0, ack => zeropad3D_CP_2152_elements(860)); -- 
    -- CP-element group 861:  transition  input  bypass 
    -- CP-element group 861: predecessors 
    -- CP-element group 861: 	859 
    -- CP-element group 861: successors 
    -- CP-element group 861: 	863 
    -- CP-element group 861:  members (1) 
      -- CP-element group 861: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/phi_stmt_1313_ack
      -- 
    phi_stmt_1313_ack_11839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 861_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1313_ack_0, ack => zeropad3D_CP_2152_elements(861)); -- 
    -- CP-element group 862:  transition  input  bypass 
    -- CP-element group 862: predecessors 
    -- CP-element group 862: 	859 
    -- CP-element group 862: successors 
    -- CP-element group 862: 	863 
    -- CP-element group 862:  members (1) 
      -- CP-element group 862: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/phi_stmt_1319_ack
      -- 
    phi_stmt_1319_ack_11840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 862_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1319_ack_0, ack => zeropad3D_CP_2152_elements(862)); -- 
    -- CP-element group 863:  join  transition  bypass 
    -- CP-element group 863: predecessors 
    -- CP-element group 863: 	860 
    -- CP-element group 863: 	861 
    -- CP-element group 863: 	862 
    -- CP-element group 863: successors 
    -- CP-element group 863: 	1 
    -- CP-element group 863:  members (1) 
      -- CP-element group 863: 	 branch_block_stmt_714/merge_stmt_1306_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_863: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_863"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(860) & zeropad3D_CP_2152_elements(861) & zeropad3D_CP_2152_elements(862);
      gj_zeropad3D_cp_element_group_863 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(863), clk => clk, reset => reset); --
    end block;
    -- CP-element group 864:  transition  input  bypass 
    -- CP-element group 864: predecessors 
    -- CP-element group 864: 	2 
    -- CP-element group 864: successors 
    -- CP-element group 864: 	866 
    -- CP-element group 864:  members (2) 
      -- CP-element group 864: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Sample/$exit
      -- CP-element group 864: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Sample/ra
      -- 
    ra_11868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 864_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_0, ack => zeropad3D_CP_2152_elements(864)); -- 
    -- CP-element group 865:  transition  input  bypass 
    -- CP-element group 865: predecessors 
    -- CP-element group 865: 	2 
    -- CP-element group 865: successors 
    -- CP-element group 865: 	866 
    -- CP-element group 865:  members (2) 
      -- CP-element group 865: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Update/$exit
      -- CP-element group 865: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/Update/ca
      -- 
    ca_11873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 865_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1468_inst_ack_1, ack => zeropad3D_CP_2152_elements(865)); -- 
    -- CP-element group 866:  join  transition  output  bypass 
    -- CP-element group 866: predecessors 
    -- CP-element group 866: 	864 
    -- CP-element group 866: 	865 
    -- CP-element group 866: successors 
    -- CP-element group 866: 	873 
    -- CP-element group 866:  members (5) 
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/$exit
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/$exit
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/$exit
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1468/SplitProtocol/$exit
      -- CP-element group 866: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_req
      -- 
    phi_stmt_1463_req_11874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1463_req_11874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(866), ack => phi_stmt_1463_req_1); -- 
    zeropad3D_cp_element_group_866: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_866"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(864) & zeropad3D_CP_2152_elements(865);
      gj_zeropad3D_cp_element_group_866 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(866), clk => clk, reset => reset); --
    end block;
    -- CP-element group 867:  transition  input  bypass 
    -- CP-element group 867: predecessors 
    -- CP-element group 867: 	2 
    -- CP-element group 867: successors 
    -- CP-element group 867: 	869 
    -- CP-element group 867:  members (2) 
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Sample/$exit
      -- CP-element group 867: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Sample/ra
      -- 
    ra_11891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 867_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1475_inst_ack_0, ack => zeropad3D_CP_2152_elements(867)); -- 
    -- CP-element group 868:  transition  input  bypass 
    -- CP-element group 868: predecessors 
    -- CP-element group 868: 	2 
    -- CP-element group 868: successors 
    -- CP-element group 868: 	869 
    -- CP-element group 868:  members (2) 
      -- CP-element group 868: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Update/$exit
      -- CP-element group 868: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/Update/ca
      -- 
    ca_11896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 868_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1475_inst_ack_1, ack => zeropad3D_CP_2152_elements(868)); -- 
    -- CP-element group 869:  join  transition  output  bypass 
    -- CP-element group 869: predecessors 
    -- CP-element group 869: 	867 
    -- CP-element group 869: 	868 
    -- CP-element group 869: successors 
    -- CP-element group 869: 	873 
    -- CP-element group 869:  members (5) 
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/$exit
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/$exit
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/$exit
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1475/SplitProtocol/$exit
      -- CP-element group 869: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_req
      -- 
    phi_stmt_1469_req_11897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1469_req_11897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(869), ack => phi_stmt_1469_req_1); -- 
    zeropad3D_cp_element_group_869: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_869"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(867) & zeropad3D_CP_2152_elements(868);
      gj_zeropad3D_cp_element_group_869 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(869), clk => clk, reset => reset); --
    end block;
    -- CP-element group 870:  transition  input  bypass 
    -- CP-element group 870: predecessors 
    -- CP-element group 870: 	2 
    -- CP-element group 870: successors 
    -- CP-element group 870: 	872 
    -- CP-element group 870:  members (2) 
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Sample/$exit
      -- CP-element group 870: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Sample/ra
      -- 
    ra_11914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 870_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1482_inst_ack_0, ack => zeropad3D_CP_2152_elements(870)); -- 
    -- CP-element group 871:  transition  input  bypass 
    -- CP-element group 871: predecessors 
    -- CP-element group 871: 	2 
    -- CP-element group 871: successors 
    -- CP-element group 871: 	872 
    -- CP-element group 871:  members (2) 
      -- CP-element group 871: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Update/$exit
      -- CP-element group 871: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/Update/ca
      -- 
    ca_11919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 871_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1482_inst_ack_1, ack => zeropad3D_CP_2152_elements(871)); -- 
    -- CP-element group 872:  join  transition  output  bypass 
    -- CP-element group 872: predecessors 
    -- CP-element group 872: 	870 
    -- CP-element group 872: 	871 
    -- CP-element group 872: successors 
    -- CP-element group 872: 	873 
    -- CP-element group 872:  members (5) 
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/$exit
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/$exit
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/$exit
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1482/SplitProtocol/$exit
      -- CP-element group 872: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_req
      -- 
    phi_stmt_1476_req_11920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1476_req_11920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(872), ack => phi_stmt_1476_req_1); -- 
    zeropad3D_cp_element_group_872: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_872"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(870) & zeropad3D_CP_2152_elements(871);
      gj_zeropad3D_cp_element_group_872 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(872), clk => clk, reset => reset); --
    end block;
    -- CP-element group 873:  join  transition  bypass 
    -- CP-element group 873: predecessors 
    -- CP-element group 873: 	866 
    -- CP-element group 873: 	869 
    -- CP-element group 873: 	872 
    -- CP-element group 873: successors 
    -- CP-element group 873: 	880 
    -- CP-element group 873:  members (1) 
      -- CP-element group 873: 	 branch_block_stmt_714/ifx_xend399_whilex_xbody244_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_873: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_873"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(866) & zeropad3D_CP_2152_elements(869) & zeropad3D_CP_2152_elements(872);
      gj_zeropad3D_cp_element_group_873 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(873), clk => clk, reset => reset); --
    end block;
    -- CP-element group 874:  transition  input  bypass 
    -- CP-element group 874: predecessors 
    -- CP-element group 874: 	153 
    -- CP-element group 874: successors 
    -- CP-element group 874: 	876 
    -- CP-element group 874:  members (2) 
      -- CP-element group 874: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Sample/$exit
      -- CP-element group 874: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Sample/ra
      -- 
    ra_11940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 874_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_0, ack => zeropad3D_CP_2152_elements(874)); -- 
    -- CP-element group 875:  transition  input  bypass 
    -- CP-element group 875: predecessors 
    -- CP-element group 875: 	153 
    -- CP-element group 875: successors 
    -- CP-element group 875: 	876 
    -- CP-element group 875:  members (2) 
      -- CP-element group 875: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Update/$exit
      -- CP-element group 875: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/Update/ca
      -- 
    ca_11945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 875_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_1, ack => zeropad3D_CP_2152_elements(875)); -- 
    -- CP-element group 876:  join  transition  output  bypass 
    -- CP-element group 876: predecessors 
    -- CP-element group 876: 	874 
    -- CP-element group 876: 	875 
    -- CP-element group 876: successors 
    -- CP-element group 876: 	879 
    -- CP-element group 876:  members (5) 
      -- CP-element group 876: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/$exit
      -- CP-element group 876: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/$exit
      -- CP-element group 876: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/$exit
      -- CP-element group 876: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_sources/type_cast_1466/SplitProtocol/$exit
      -- CP-element group 876: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1463/phi_stmt_1463_req
      -- 
    phi_stmt_1463_req_11946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1463_req_11946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(876), ack => phi_stmt_1463_req_0); -- 
    zeropad3D_cp_element_group_876: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_876"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(874) & zeropad3D_CP_2152_elements(875);
      gj_zeropad3D_cp_element_group_876 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(876), clk => clk, reset => reset); --
    end block;
    -- CP-element group 877:  transition  output  delay-element  bypass 
    -- CP-element group 877: predecessors 
    -- CP-element group 877: 	153 
    -- CP-element group 877: successors 
    -- CP-element group 877: 	879 
    -- CP-element group 877:  members (4) 
      -- CP-element group 877: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1469/$exit
      -- CP-element group 877: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/$exit
      -- CP-element group 877: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_sources/type_cast_1473_konst_delay_trans
      -- CP-element group 877: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1469/phi_stmt_1469_req
      -- 
    phi_stmt_1469_req_11954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1469_req_11954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(877), ack => phi_stmt_1469_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(877) is a control-delay.
    cp_element_877_delay: control_delay_element  generic map(name => " 877_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(153), ack => zeropad3D_CP_2152_elements(877), clk => clk, reset =>reset);
    -- CP-element group 878:  transition  output  delay-element  bypass 
    -- CP-element group 878: predecessors 
    -- CP-element group 878: 	153 
    -- CP-element group 878: successors 
    -- CP-element group 878: 	879 
    -- CP-element group 878:  members (4) 
      -- CP-element group 878: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1476/$exit
      -- CP-element group 878: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/$exit
      -- CP-element group 878: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_sources/type_cast_1480_konst_delay_trans
      -- CP-element group 878: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/phi_stmt_1476/phi_stmt_1476_req
      -- 
    phi_stmt_1476_req_11962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1476_req_11962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(878), ack => phi_stmt_1476_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(878) is a control-delay.
    cp_element_878_delay: control_delay_element  generic map(name => " 878_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(153), ack => zeropad3D_CP_2152_elements(878), clk => clk, reset =>reset);
    -- CP-element group 879:  join  transition  bypass 
    -- CP-element group 879: predecessors 
    -- CP-element group 879: 	876 
    -- CP-element group 879: 	877 
    -- CP-element group 879: 	878 
    -- CP-element group 879: successors 
    -- CP-element group 879: 	880 
    -- CP-element group 879:  members (1) 
      -- CP-element group 879: 	 branch_block_stmt_714/whilex_xend_whilex_xbody244_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_879: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_879"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(876) & zeropad3D_CP_2152_elements(877) & zeropad3D_CP_2152_elements(878);
      gj_zeropad3D_cp_element_group_879 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(879), clk => clk, reset => reset); --
    end block;
    -- CP-element group 880:  merge  fork  transition  place  bypass 
    -- CP-element group 880: predecessors 
    -- CP-element group 880: 	873 
    -- CP-element group 880: 	879 
    -- CP-element group 880: successors 
    -- CP-element group 880: 	881 
    -- CP-element group 880: 	882 
    -- CP-element group 880: 	883 
    -- CP-element group 880:  members (2) 
      -- CP-element group 880: 	 branch_block_stmt_714/merge_stmt_1462_PhiReqMerge
      -- CP-element group 880: 	 branch_block_stmt_714/merge_stmt_1462_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(880) <= OrReduce(zeropad3D_CP_2152_elements(873) & zeropad3D_CP_2152_elements(879));
    -- CP-element group 881:  transition  input  bypass 
    -- CP-element group 881: predecessors 
    -- CP-element group 881: 	880 
    -- CP-element group 881: successors 
    -- CP-element group 881: 	884 
    -- CP-element group 881:  members (1) 
      -- CP-element group 881: 	 branch_block_stmt_714/merge_stmt_1462_PhiAck/phi_stmt_1463_ack
      -- 
    phi_stmt_1463_ack_11967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 881_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1463_ack_0, ack => zeropad3D_CP_2152_elements(881)); -- 
    -- CP-element group 882:  transition  input  bypass 
    -- CP-element group 882: predecessors 
    -- CP-element group 882: 	880 
    -- CP-element group 882: successors 
    -- CP-element group 882: 	884 
    -- CP-element group 882:  members (1) 
      -- CP-element group 882: 	 branch_block_stmt_714/merge_stmt_1462_PhiAck/phi_stmt_1469_ack
      -- 
    phi_stmt_1469_ack_11968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 882_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1469_ack_0, ack => zeropad3D_CP_2152_elements(882)); -- 
    -- CP-element group 883:  transition  input  bypass 
    -- CP-element group 883: predecessors 
    -- CP-element group 883: 	880 
    -- CP-element group 883: successors 
    -- CP-element group 883: 	884 
    -- CP-element group 883:  members (1) 
      -- CP-element group 883: 	 branch_block_stmt_714/merge_stmt_1462_PhiAck/phi_stmt_1476_ack
      -- 
    phi_stmt_1476_ack_11969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 883_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1476_ack_0, ack => zeropad3D_CP_2152_elements(883)); -- 
    -- CP-element group 884:  join  fork  transition  place  output  bypass 
    -- CP-element group 884: predecessors 
    -- CP-element group 884: 	881 
    -- CP-element group 884: 	882 
    -- CP-element group 884: 	883 
    -- CP-element group 884: successors 
    -- CP-element group 884: 	154 
    -- CP-element group 884: 	155 
    -- CP-element group 884:  members (10) 
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495__entry__
      -- CP-element group 884: 	 branch_block_stmt_714/merge_stmt_1462__exit__
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/$entry
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_sample_start_
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_update_start_
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Sample/$entry
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Sample/rr
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Update/$entry
      -- CP-element group 884: 	 branch_block_stmt_714/assign_stmt_1488_to_assign_stmt_1495/type_cast_1487_Update/cr
      -- CP-element group 884: 	 branch_block_stmt_714/merge_stmt_1462_PhiAck/$exit
      -- 
    rr_4209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(884), ack => type_cast_1487_inst_req_0); -- 
    cr_4214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(884), ack => type_cast_1487_inst_req_1); -- 
    zeropad3D_cp_element_group_884: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_884"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(881) & zeropad3D_CP_2152_elements(882) & zeropad3D_CP_2152_elements(883);
      gj_zeropad3D_cp_element_group_884 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(884), clk => clk, reset => reset); --
    end block;
    -- CP-element group 885:  merge  fork  transition  place  output  bypass 
    -- CP-element group 885: predecessors 
    -- CP-element group 885: 	156 
    -- CP-element group 885: 	163 
    -- CP-element group 885: 	166 
    -- CP-element group 885: 	173 
    -- CP-element group 885: successors 
    -- CP-element group 885: 	174 
    -- CP-element group 885: 	175 
    -- CP-element group 885: 	176 
    -- CP-element group 885: 	177 
    -- CP-element group 885: 	180 
    -- CP-element group 885: 	182 
    -- CP-element group 885: 	184 
    -- CP-element group 885: 	186 
    -- CP-element group 885:  members (33) 
      -- CP-element group 885: 	 branch_block_stmt_714/merge_stmt_1579__exit__
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635__entry__
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Update/req
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_sample_start_
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_Update/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_update_start_
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/array_obj_ref_1628_final_index_sum_regn_update_start
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/word_access_complete/word_0/cr
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/word_access_complete/word_0/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/word_access_complete/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/ptr_deref_1632_Update/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_complete/req
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_complete/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/addr_of_1629_update_start_
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Update/cr
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_Update/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1622_update_start_
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Update/cr
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Update/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Sample/rr
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_Sample/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_update_start_
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1588_sample_start_
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Update/cr
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Update/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Sample/rr
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_Sample/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/assign_stmt_1584_to_assign_stmt_1635/type_cast_1583_update_start_
      -- CP-element group 885: 	 branch_block_stmt_714/merge_stmt_1579_PhiReqMerge
      -- CP-element group 885: 	 branch_block_stmt_714/merge_stmt_1579_PhiAck/$entry
      -- CP-element group 885: 	 branch_block_stmt_714/merge_stmt_1579_PhiAck/$exit
      -- CP-element group 885: 	 branch_block_stmt_714/merge_stmt_1579_PhiAck/dummy
      -- 
    req_4483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => array_obj_ref_1628_index_offset_req_1); -- 
    cr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => ptr_deref_1632_store_0_req_1); -- 
    req_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => addr_of_1629_final_reg_req_1); -- 
    cr_4452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => type_cast_1622_inst_req_1); -- 
    cr_4438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => type_cast_1588_inst_req_1); -- 
    rr_4433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => type_cast_1588_inst_req_0); -- 
    cr_4424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => type_cast_1583_inst_req_1); -- 
    rr_4419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(885), ack => type_cast_1583_inst_req_0); -- 
    zeropad3D_CP_2152_elements(885) <= OrReduce(zeropad3D_CP_2152_elements(156) & zeropad3D_CP_2152_elements(163) & zeropad3D_CP_2152_elements(166) & zeropad3D_CP_2152_elements(173));
    -- CP-element group 886:  merge  fork  transition  place  output  bypass 
    -- CP-element group 886: predecessors 
    -- CP-element group 886: 	187 
    -- CP-element group 886: 	207 
    -- CP-element group 886: successors 
    -- CP-element group 886: 	208 
    -- CP-element group 886: 	209 
    -- CP-element group 886:  members (13) 
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762__entry__
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1744__exit__
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/$entry
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_sample_start_
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_update_start_
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Sample/$entry
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Sample/rr
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Update/$entry
      -- CP-element group 886: 	 branch_block_stmt_714/assign_stmt_1749_to_assign_stmt_1762/type_cast_1748_Update/cr
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1744_PhiReqMerge
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1744_PhiAck/$entry
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1744_PhiAck/$exit
      -- CP-element group 886: 	 branch_block_stmt_714/merge_stmt_1744_PhiAck/dummy
      -- 
    rr_4797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(886), ack => type_cast_1748_inst_req_0); -- 
    cr_4802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(886), ack => type_cast_1748_inst_req_1); -- 
    zeropad3D_CP_2152_elements(886) <= OrReduce(zeropad3D_CP_2152_elements(187) & zeropad3D_CP_2152_elements(207));
    -- CP-element group 887:  transition  output  delay-element  bypass 
    -- CP-element group 887: predecessors 
    -- CP-element group 887: 	229 
    -- CP-element group 887: successors 
    -- CP-element group 887: 	894 
    -- CP-element group 887:  members (4) 
      -- CP-element group 887: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1868/$exit
      -- CP-element group 887: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$exit
      -- CP-element group 887: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1874_konst_delay_trans
      -- CP-element group 887: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_req
      -- 
    phi_stmt_1868_req_12080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_req_12080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(887), ack => phi_stmt_1868_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(887) is a control-delay.
    cp_element_887_delay: control_delay_element  generic map(name => " 887_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(229), ack => zeropad3D_CP_2152_elements(887), clk => clk, reset =>reset);
    -- CP-element group 888:  transition  input  bypass 
    -- CP-element group 888: predecessors 
    -- CP-element group 888: 	229 
    -- CP-element group 888: successors 
    -- CP-element group 888: 	890 
    -- CP-element group 888:  members (2) 
      -- CP-element group 888: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Sample/$exit
      -- CP-element group 888: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Sample/ra
      -- 
    ra_12097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 888_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_0, ack => zeropad3D_CP_2152_elements(888)); -- 
    -- CP-element group 889:  transition  input  bypass 
    -- CP-element group 889: predecessors 
    -- CP-element group 889: 	229 
    -- CP-element group 889: successors 
    -- CP-element group 889: 	890 
    -- CP-element group 889:  members (2) 
      -- CP-element group 889: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Update/$exit
      -- CP-element group 889: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/Update/ca
      -- 
    ca_12102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 889_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_1, ack => zeropad3D_CP_2152_elements(889)); -- 
    -- CP-element group 890:  join  transition  output  bypass 
    -- CP-element group 890: predecessors 
    -- CP-element group 890: 	888 
    -- CP-element group 890: 	889 
    -- CP-element group 890: successors 
    -- CP-element group 890: 	894 
    -- CP-element group 890:  members (5) 
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/$exit
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$exit
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/$exit
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1867/SplitProtocol/$exit
      -- CP-element group 890: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_req
      -- 
    phi_stmt_1862_req_12103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1862_req_12103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(890), ack => phi_stmt_1862_req_1); -- 
    zeropad3D_cp_element_group_890: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_890"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(888) & zeropad3D_CP_2152_elements(889);
      gj_zeropad3D_cp_element_group_890 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(890), clk => clk, reset => reset); --
    end block;
    -- CP-element group 891:  transition  input  bypass 
    -- CP-element group 891: predecessors 
    -- CP-element group 891: 	229 
    -- CP-element group 891: successors 
    -- CP-element group 891: 	893 
    -- CP-element group 891:  members (2) 
      -- CP-element group 891: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Sample/$exit
      -- CP-element group 891: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Sample/ra
      -- 
    ra_12120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 891_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1861_inst_ack_0, ack => zeropad3D_CP_2152_elements(891)); -- 
    -- CP-element group 892:  transition  input  bypass 
    -- CP-element group 892: predecessors 
    -- CP-element group 892: 	229 
    -- CP-element group 892: successors 
    -- CP-element group 892: 	893 
    -- CP-element group 892:  members (2) 
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Update/$exit
      -- CP-element group 892: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/Update/ca
      -- 
    ca_12125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 892_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1861_inst_ack_1, ack => zeropad3D_CP_2152_elements(892)); -- 
    -- CP-element group 893:  join  transition  output  bypass 
    -- CP-element group 893: predecessors 
    -- CP-element group 893: 	891 
    -- CP-element group 893: 	892 
    -- CP-element group 893: successors 
    -- CP-element group 893: 	894 
    -- CP-element group 893:  members (5) 
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/$exit
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/$exit
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/$exit
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1861/SplitProtocol/$exit
      -- CP-element group 893: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_req
      -- 
    phi_stmt_1856_req_12126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1856_req_12126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(893), ack => phi_stmt_1856_req_1); -- 
    zeropad3D_cp_element_group_893: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_893"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(891) & zeropad3D_CP_2152_elements(892);
      gj_zeropad3D_cp_element_group_893 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(893), clk => clk, reset => reset); --
    end block;
    -- CP-element group 894:  join  transition  bypass 
    -- CP-element group 894: predecessors 
    -- CP-element group 894: 	887 
    -- CP-element group 894: 	890 
    -- CP-element group 894: 	893 
    -- CP-element group 894: successors 
    -- CP-element group 894: 	905 
    -- CP-element group 894:  members (1) 
      -- CP-element group 894: 	 branch_block_stmt_714/ifx_xelse363_ifx_xend399_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_894: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_894"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(887) & zeropad3D_CP_2152_elements(890) & zeropad3D_CP_2152_elements(893);
      gj_zeropad3D_cp_element_group_894 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(894), clk => clk, reset => reset); --
    end block;
    -- CP-element group 895:  transition  input  bypass 
    -- CP-element group 895: predecessors 
    -- CP-element group 895: 	210 
    -- CP-element group 895: successors 
    -- CP-element group 895: 	897 
    -- CP-element group 895:  members (2) 
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Sample/$exit
      -- CP-element group 895: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Sample/ra
      -- 
    ra_12146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 895_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1871_inst_ack_0, ack => zeropad3D_CP_2152_elements(895)); -- 
    -- CP-element group 896:  transition  input  bypass 
    -- CP-element group 896: predecessors 
    -- CP-element group 896: 	210 
    -- CP-element group 896: successors 
    -- CP-element group 896: 	897 
    -- CP-element group 896:  members (2) 
      -- CP-element group 896: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Update/$exit
      -- CP-element group 896: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/Update/ca
      -- 
    ca_12151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 896_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1871_inst_ack_1, ack => zeropad3D_CP_2152_elements(896)); -- 
    -- CP-element group 897:  join  transition  output  bypass 
    -- CP-element group 897: predecessors 
    -- CP-element group 897: 	895 
    -- CP-element group 897: 	896 
    -- CP-element group 897: successors 
    -- CP-element group 897: 	904 
    -- CP-element group 897:  members (5) 
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/$exit
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/$exit
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/$exit
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_sources/type_cast_1871/SplitProtocol/$exit
      -- CP-element group 897: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1868/phi_stmt_1868_req
      -- 
    phi_stmt_1868_req_12152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_req_12152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(897), ack => phi_stmt_1868_req_0); -- 
    zeropad3D_cp_element_group_897: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_897"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(895) & zeropad3D_CP_2152_elements(896);
      gj_zeropad3D_cp_element_group_897 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(897), clk => clk, reset => reset); --
    end block;
    -- CP-element group 898:  transition  input  bypass 
    -- CP-element group 898: predecessors 
    -- CP-element group 898: 	210 
    -- CP-element group 898: successors 
    -- CP-element group 898: 	900 
    -- CP-element group 898:  members (2) 
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Sample/$exit
      -- CP-element group 898: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Sample/ra
      -- 
    ra_12169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 898_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_0, ack => zeropad3D_CP_2152_elements(898)); -- 
    -- CP-element group 899:  transition  input  bypass 
    -- CP-element group 899: predecessors 
    -- CP-element group 899: 	210 
    -- CP-element group 899: successors 
    -- CP-element group 899: 	900 
    -- CP-element group 899:  members (2) 
      -- CP-element group 899: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Update/$exit
      -- CP-element group 899: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/Update/ca
      -- 
    ca_12174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 899_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_1, ack => zeropad3D_CP_2152_elements(899)); -- 
    -- CP-element group 900:  join  transition  output  bypass 
    -- CP-element group 900: predecessors 
    -- CP-element group 900: 	898 
    -- CP-element group 900: 	899 
    -- CP-element group 900: successors 
    -- CP-element group 900: 	904 
    -- CP-element group 900:  members (5) 
      -- CP-element group 900: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/$exit
      -- CP-element group 900: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$exit
      -- CP-element group 900: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/$exit
      -- CP-element group 900: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1865/SplitProtocol/$exit
      -- CP-element group 900: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1862/phi_stmt_1862_req
      -- 
    phi_stmt_1862_req_12175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1862_req_12175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(900), ack => phi_stmt_1862_req_0); -- 
    zeropad3D_cp_element_group_900: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_900"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(898) & zeropad3D_CP_2152_elements(899);
      gj_zeropad3D_cp_element_group_900 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(900), clk => clk, reset => reset); --
    end block;
    -- CP-element group 901:  transition  input  bypass 
    -- CP-element group 901: predecessors 
    -- CP-element group 901: 	210 
    -- CP-element group 901: successors 
    -- CP-element group 901: 	903 
    -- CP-element group 901:  members (2) 
      -- CP-element group 901: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Sample/$exit
      -- CP-element group 901: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Sample/ra
      -- 
    ra_12192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 901_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1859_inst_ack_0, ack => zeropad3D_CP_2152_elements(901)); -- 
    -- CP-element group 902:  transition  input  bypass 
    -- CP-element group 902: predecessors 
    -- CP-element group 902: 	210 
    -- CP-element group 902: successors 
    -- CP-element group 902: 	903 
    -- CP-element group 902:  members (2) 
      -- CP-element group 902: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Update/$exit
      -- CP-element group 902: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/Update/ca
      -- 
    ca_12197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 902_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1859_inst_ack_1, ack => zeropad3D_CP_2152_elements(902)); -- 
    -- CP-element group 903:  join  transition  output  bypass 
    -- CP-element group 903: predecessors 
    -- CP-element group 903: 	901 
    -- CP-element group 903: 	902 
    -- CP-element group 903: successors 
    -- CP-element group 903: 	904 
    -- CP-element group 903:  members (5) 
      -- CP-element group 903: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/$exit
      -- CP-element group 903: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/$exit
      -- CP-element group 903: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/$exit
      -- CP-element group 903: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_sources/type_cast_1859/SplitProtocol/$exit
      -- CP-element group 903: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/phi_stmt_1856/phi_stmt_1856_req
      -- 
    phi_stmt_1856_req_12198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1856_req_12198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(903), ack => phi_stmt_1856_req_0); -- 
    zeropad3D_cp_element_group_903: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_903"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(901) & zeropad3D_CP_2152_elements(902);
      gj_zeropad3D_cp_element_group_903 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(903), clk => clk, reset => reset); --
    end block;
    -- CP-element group 904:  join  transition  bypass 
    -- CP-element group 904: predecessors 
    -- CP-element group 904: 	897 
    -- CP-element group 904: 	900 
    -- CP-element group 904: 	903 
    -- CP-element group 904: successors 
    -- CP-element group 904: 	905 
    -- CP-element group 904:  members (1) 
      -- CP-element group 904: 	 branch_block_stmt_714/ifx_xthen358_ifx_xend399_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_904: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_904"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(897) & zeropad3D_CP_2152_elements(900) & zeropad3D_CP_2152_elements(903);
      gj_zeropad3D_cp_element_group_904 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(904), clk => clk, reset => reset); --
    end block;
    -- CP-element group 905:  merge  fork  transition  place  bypass 
    -- CP-element group 905: predecessors 
    -- CP-element group 905: 	894 
    -- CP-element group 905: 	904 
    -- CP-element group 905: successors 
    -- CP-element group 905: 	906 
    -- CP-element group 905: 	907 
    -- CP-element group 905: 	908 
    -- CP-element group 905:  members (2) 
      -- CP-element group 905: 	 branch_block_stmt_714/merge_stmt_1855_PhiReqMerge
      -- CP-element group 905: 	 branch_block_stmt_714/merge_stmt_1855_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(905) <= OrReduce(zeropad3D_CP_2152_elements(894) & zeropad3D_CP_2152_elements(904));
    -- CP-element group 906:  transition  input  bypass 
    -- CP-element group 906: predecessors 
    -- CP-element group 906: 	905 
    -- CP-element group 906: successors 
    -- CP-element group 906: 	909 
    -- CP-element group 906:  members (1) 
      -- CP-element group 906: 	 branch_block_stmt_714/merge_stmt_1855_PhiAck/phi_stmt_1856_ack
      -- 
    phi_stmt_1856_ack_12203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 906_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1856_ack_0, ack => zeropad3D_CP_2152_elements(906)); -- 
    -- CP-element group 907:  transition  input  bypass 
    -- CP-element group 907: predecessors 
    -- CP-element group 907: 	905 
    -- CP-element group 907: successors 
    -- CP-element group 907: 	909 
    -- CP-element group 907:  members (1) 
      -- CP-element group 907: 	 branch_block_stmt_714/merge_stmt_1855_PhiAck/phi_stmt_1862_ack
      -- 
    phi_stmt_1862_ack_12204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 907_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1862_ack_0, ack => zeropad3D_CP_2152_elements(907)); -- 
    -- CP-element group 908:  transition  input  bypass 
    -- CP-element group 908: predecessors 
    -- CP-element group 908: 	905 
    -- CP-element group 908: successors 
    -- CP-element group 908: 	909 
    -- CP-element group 908:  members (1) 
      -- CP-element group 908: 	 branch_block_stmt_714/merge_stmt_1855_PhiAck/phi_stmt_1868_ack
      -- 
    phi_stmt_1868_ack_12205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 908_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1868_ack_0, ack => zeropad3D_CP_2152_elements(908)); -- 
    -- CP-element group 909:  join  transition  bypass 
    -- CP-element group 909: predecessors 
    -- CP-element group 909: 	906 
    -- CP-element group 909: 	907 
    -- CP-element group 909: 	908 
    -- CP-element group 909: successors 
    -- CP-element group 909: 	2 
    -- CP-element group 909:  members (1) 
      -- CP-element group 909: 	 branch_block_stmt_714/merge_stmt_1855_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_909: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_909"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(906) & zeropad3D_CP_2152_elements(907) & zeropad3D_CP_2152_elements(908);
      gj_zeropad3D_cp_element_group_909 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(909), clk => clk, reset => reset); --
    end block;
    -- CP-element group 910:  transition  input  bypass 
    -- CP-element group 910: predecessors 
    -- CP-element group 910: 	3 
    -- CP-element group 910: successors 
    -- CP-element group 910: 	912 
    -- CP-element group 910:  members (2) 
      -- CP-element group 910: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Sample/$exit
      -- CP-element group 910: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Sample/ra
      -- 
    ra_12233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 910_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_0, ack => zeropad3D_CP_2152_elements(910)); -- 
    -- CP-element group 911:  transition  input  bypass 
    -- CP-element group 911: predecessors 
    -- CP-element group 911: 	3 
    -- CP-element group 911: successors 
    -- CP-element group 911: 	912 
    -- CP-element group 911:  members (2) 
      -- CP-element group 911: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Update/$exit
      -- CP-element group 911: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/Update/ca
      -- 
    ca_12238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 911_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_1, ack => zeropad3D_CP_2152_elements(911)); -- 
    -- CP-element group 912:  join  transition  output  bypass 
    -- CP-element group 912: predecessors 
    -- CP-element group 912: 	910 
    -- CP-element group 912: 	911 
    -- CP-element group 912: successors 
    -- CP-element group 912: 	919 
    -- CP-element group 912:  members (5) 
      -- CP-element group 912: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/$exit
      -- CP-element group 912: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/$exit
      -- CP-element group 912: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/$exit
      -- CP-element group 912: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2018/SplitProtocol/$exit
      -- CP-element group 912: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_req
      -- 
    phi_stmt_2015_req_12239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2015_req_12239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(912), ack => phi_stmt_2015_req_0); -- 
    zeropad3D_cp_element_group_912: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_912"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(910) & zeropad3D_CP_2152_elements(911);
      gj_zeropad3D_cp_element_group_912 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(912), clk => clk, reset => reset); --
    end block;
    -- CP-element group 913:  transition  input  bypass 
    -- CP-element group 913: predecessors 
    -- CP-element group 913: 	3 
    -- CP-element group 913: successors 
    -- CP-element group 913: 	915 
    -- CP-element group 913:  members (2) 
      -- CP-element group 913: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Sample/$exit
      -- CP-element group 913: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Sample/ra
      -- 
    ra_12256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 913_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_0, ack => zeropad3D_CP_2152_elements(913)); -- 
    -- CP-element group 914:  transition  input  bypass 
    -- CP-element group 914: predecessors 
    -- CP-element group 914: 	3 
    -- CP-element group 914: successors 
    -- CP-element group 914: 	915 
    -- CP-element group 914:  members (2) 
      -- CP-element group 914: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Update/$exit
      -- CP-element group 914: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/Update/ca
      -- 
    ca_12261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 914_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_1, ack => zeropad3D_CP_2152_elements(914)); -- 
    -- CP-element group 915:  join  transition  output  bypass 
    -- CP-element group 915: predecessors 
    -- CP-element group 915: 	913 
    -- CP-element group 915: 	914 
    -- CP-element group 915: successors 
    -- CP-element group 915: 	919 
    -- CP-element group 915:  members (5) 
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/$exit
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/$exit
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/$exit
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2031/SplitProtocol/$exit
      -- CP-element group 915: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_req
      -- 
    phi_stmt_2028_req_12262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2028_req_12262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(915), ack => phi_stmt_2028_req_0); -- 
    zeropad3D_cp_element_group_915: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_915"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(913) & zeropad3D_CP_2152_elements(914);
      gj_zeropad3D_cp_element_group_915 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(915), clk => clk, reset => reset); --
    end block;
    -- CP-element group 916:  transition  input  bypass 
    -- CP-element group 916: predecessors 
    -- CP-element group 916: 	3 
    -- CP-element group 916: successors 
    -- CP-element group 916: 	918 
    -- CP-element group 916:  members (2) 
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Sample/$exit
      -- CP-element group 916: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Sample/ra
      -- 
    ra_12279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 916_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2027_inst_ack_0, ack => zeropad3D_CP_2152_elements(916)); -- 
    -- CP-element group 917:  transition  input  bypass 
    -- CP-element group 917: predecessors 
    -- CP-element group 917: 	3 
    -- CP-element group 917: successors 
    -- CP-element group 917: 	918 
    -- CP-element group 917:  members (2) 
      -- CP-element group 917: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Update/$exit
      -- CP-element group 917: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/Update/ca
      -- 
    ca_12284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 917_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2027_inst_ack_1, ack => zeropad3D_CP_2152_elements(917)); -- 
    -- CP-element group 918:  join  transition  output  bypass 
    -- CP-element group 918: predecessors 
    -- CP-element group 918: 	916 
    -- CP-element group 918: 	917 
    -- CP-element group 918: successors 
    -- CP-element group 918: 	919 
    -- CP-element group 918:  members (5) 
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/$exit
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/$exit
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/$exit
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2027/SplitProtocol/$exit
      -- CP-element group 918: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_req
      -- 
    phi_stmt_2022_req_12285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2022_req_12285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(918), ack => phi_stmt_2022_req_1); -- 
    zeropad3D_cp_element_group_918: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_918"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(916) & zeropad3D_CP_2152_elements(917);
      gj_zeropad3D_cp_element_group_918 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(918), clk => clk, reset => reset); --
    end block;
    -- CP-element group 919:  join  transition  bypass 
    -- CP-element group 919: predecessors 
    -- CP-element group 919: 	912 
    -- CP-element group 919: 	915 
    -- CP-element group 919: 	918 
    -- CP-element group 919: successors 
    -- CP-element group 919: 	926 
    -- CP-element group 919:  members (1) 
      -- CP-element group 919: 	 branch_block_stmt_714/ifx_xend617_whilex_xbody460_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_919: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_919"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(912) & zeropad3D_CP_2152_elements(915) & zeropad3D_CP_2152_elements(918);
      gj_zeropad3D_cp_element_group_919 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(919), clk => clk, reset => reset); --
    end block;
    -- CP-element group 920:  transition  output  delay-element  bypass 
    -- CP-element group 920: predecessors 
    -- CP-element group 920: 	250 
    -- CP-element group 920: successors 
    -- CP-element group 920: 	925 
    -- CP-element group 920:  members (4) 
      -- CP-element group 920: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2015/$exit
      -- CP-element group 920: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/$exit
      -- CP-element group 920: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_sources/type_cast_2021_konst_delay_trans
      -- CP-element group 920: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2015/phi_stmt_2015_req
      -- 
    phi_stmt_2015_req_12296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2015_req_12296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(920), ack => phi_stmt_2015_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(920) is a control-delay.
    cp_element_920_delay: control_delay_element  generic map(name => " 920_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(250), ack => zeropad3D_CP_2152_elements(920), clk => clk, reset =>reset);
    -- CP-element group 921:  transition  output  delay-element  bypass 
    -- CP-element group 921: predecessors 
    -- CP-element group 921: 	250 
    -- CP-element group 921: successors 
    -- CP-element group 921: 	925 
    -- CP-element group 921:  members (4) 
      -- CP-element group 921: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2028/$exit
      -- CP-element group 921: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/$exit
      -- CP-element group 921: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_sources/type_cast_2034_konst_delay_trans
      -- CP-element group 921: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2028/phi_stmt_2028_req
      -- 
    phi_stmt_2028_req_12304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2028_req_12304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(921), ack => phi_stmt_2028_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(921) is a control-delay.
    cp_element_921_delay: control_delay_element  generic map(name => " 921_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(250), ack => zeropad3D_CP_2152_elements(921), clk => clk, reset =>reset);
    -- CP-element group 922:  transition  input  bypass 
    -- CP-element group 922: predecessors 
    -- CP-element group 922: 	250 
    -- CP-element group 922: successors 
    -- CP-element group 922: 	924 
    -- CP-element group 922:  members (2) 
      -- CP-element group 922: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Sample/$exit
      -- CP-element group 922: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Sample/ra
      -- 
    ra_12321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 922_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_0, ack => zeropad3D_CP_2152_elements(922)); -- 
    -- CP-element group 923:  transition  input  bypass 
    -- CP-element group 923: predecessors 
    -- CP-element group 923: 	250 
    -- CP-element group 923: successors 
    -- CP-element group 923: 	924 
    -- CP-element group 923:  members (2) 
      -- CP-element group 923: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Update/$exit
      -- CP-element group 923: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/Update/ca
      -- 
    ca_12326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 923_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_1, ack => zeropad3D_CP_2152_elements(923)); -- 
    -- CP-element group 924:  join  transition  output  bypass 
    -- CP-element group 924: predecessors 
    -- CP-element group 924: 	922 
    -- CP-element group 924: 	923 
    -- CP-element group 924: successors 
    -- CP-element group 924: 	925 
    -- CP-element group 924:  members (5) 
      -- CP-element group 924: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/$exit
      -- CP-element group 924: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/$exit
      -- CP-element group 924: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/$exit
      -- CP-element group 924: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_sources/type_cast_2025/SplitProtocol/$exit
      -- CP-element group 924: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/phi_stmt_2022/phi_stmt_2022_req
      -- 
    phi_stmt_2022_req_12327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2022_req_12327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(924), ack => phi_stmt_2022_req_0); -- 
    zeropad3D_cp_element_group_924: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_924"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(922) & zeropad3D_CP_2152_elements(923);
      gj_zeropad3D_cp_element_group_924 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(924), clk => clk, reset => reset); --
    end block;
    -- CP-element group 925:  join  transition  bypass 
    -- CP-element group 925: predecessors 
    -- CP-element group 925: 	920 
    -- CP-element group 925: 	921 
    -- CP-element group 925: 	924 
    -- CP-element group 925: successors 
    -- CP-element group 925: 	926 
    -- CP-element group 925:  members (1) 
      -- CP-element group 925: 	 branch_block_stmt_714/whilex_xend400_whilex_xbody460_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_925: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_925"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(920) & zeropad3D_CP_2152_elements(921) & zeropad3D_CP_2152_elements(924);
      gj_zeropad3D_cp_element_group_925 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(925), clk => clk, reset => reset); --
    end block;
    -- CP-element group 926:  merge  fork  transition  place  bypass 
    -- CP-element group 926: predecessors 
    -- CP-element group 926: 	919 
    -- CP-element group 926: 	925 
    -- CP-element group 926: successors 
    -- CP-element group 926: 	927 
    -- CP-element group 926: 	928 
    -- CP-element group 926: 	929 
    -- CP-element group 926:  members (2) 
      -- CP-element group 926: 	 branch_block_stmt_714/merge_stmt_2014_PhiReqMerge
      -- CP-element group 926: 	 branch_block_stmt_714/merge_stmt_2014_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(926) <= OrReduce(zeropad3D_CP_2152_elements(919) & zeropad3D_CP_2152_elements(925));
    -- CP-element group 927:  transition  input  bypass 
    -- CP-element group 927: predecessors 
    -- CP-element group 927: 	926 
    -- CP-element group 927: successors 
    -- CP-element group 927: 	930 
    -- CP-element group 927:  members (1) 
      -- CP-element group 927: 	 branch_block_stmt_714/merge_stmt_2014_PhiAck/phi_stmt_2015_ack
      -- 
    phi_stmt_2015_ack_12332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 927_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2015_ack_0, ack => zeropad3D_CP_2152_elements(927)); -- 
    -- CP-element group 928:  transition  input  bypass 
    -- CP-element group 928: predecessors 
    -- CP-element group 928: 	926 
    -- CP-element group 928: successors 
    -- CP-element group 928: 	930 
    -- CP-element group 928:  members (1) 
      -- CP-element group 928: 	 branch_block_stmt_714/merge_stmt_2014_PhiAck/phi_stmt_2022_ack
      -- 
    phi_stmt_2022_ack_12333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 928_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2022_ack_0, ack => zeropad3D_CP_2152_elements(928)); -- 
    -- CP-element group 929:  transition  input  bypass 
    -- CP-element group 929: predecessors 
    -- CP-element group 929: 	926 
    -- CP-element group 929: successors 
    -- CP-element group 929: 	930 
    -- CP-element group 929:  members (1) 
      -- CP-element group 929: 	 branch_block_stmt_714/merge_stmt_2014_PhiAck/phi_stmt_2028_ack
      -- 
    phi_stmt_2028_ack_12334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 929_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2028_ack_0, ack => zeropad3D_CP_2152_elements(929)); -- 
    -- CP-element group 930:  join  fork  transition  place  output  bypass 
    -- CP-element group 930: predecessors 
    -- CP-element group 930: 	927 
    -- CP-element group 930: 	928 
    -- CP-element group 930: 	929 
    -- CP-element group 930: successors 
    -- CP-element group 930: 	251 
    -- CP-element group 930: 	252 
    -- CP-element group 930:  members (10) 
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047__entry__
      -- CP-element group 930: 	 branch_block_stmt_714/merge_stmt_2014__exit__
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/$entry
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_sample_start_
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_update_start_
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Sample/$entry
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Sample/rr
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Update/$entry
      -- CP-element group 930: 	 branch_block_stmt_714/assign_stmt_2040_to_assign_stmt_2047/type_cast_2039_Update/cr
      -- CP-element group 930: 	 branch_block_stmt_714/merge_stmt_2014_PhiAck/$exit
      -- 
    rr_5285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(930), ack => type_cast_2039_inst_req_0); -- 
    cr_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(930), ack => type_cast_2039_inst_req_1); -- 
    zeropad3D_cp_element_group_930: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_930"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(927) & zeropad3D_CP_2152_elements(928) & zeropad3D_CP_2152_elements(929);
      gj_zeropad3D_cp_element_group_930 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(930), clk => clk, reset => reset); --
    end block;
    -- CP-element group 931:  merge  fork  transition  place  output  bypass 
    -- CP-element group 931: predecessors 
    -- CP-element group 931: 	253 
    -- CP-element group 931: 	260 
    -- CP-element group 931: 	263 
    -- CP-element group 931: 	270 
    -- CP-element group 931: successors 
    -- CP-element group 931: 	272 
    -- CP-element group 931: 	273 
    -- CP-element group 931: 	274 
    -- CP-element group 931: 	283 
    -- CP-element group 931: 	271 
    -- CP-element group 931: 	277 
    -- CP-element group 931: 	279 
    -- CP-element group 931: 	281 
    -- CP-element group 931:  members (33) 
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193__entry__
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2137__exit__
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Sample/rr
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Update/cr
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Update/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/word_access_complete/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Sample/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Update/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Sample/rr
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_Sample/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_update_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_update_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2146_sample_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Update/cr
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/word_access_complete/word_0/cr
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_update_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_complete/req
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/ptr_deref_2190_Update/word_access_complete/word_0/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_complete/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_sample_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/addr_of_2187_update_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Update/req
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_Update/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_Update/cr
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/array_obj_ref_2186_final_index_sum_regn_update_start
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2180_update_start_
      -- CP-element group 931: 	 branch_block_stmt_714/assign_stmt_2142_to_assign_stmt_2193/type_cast_2141_Update/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2137_PhiReqMerge
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2137_PhiAck/$entry
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2137_PhiAck/$exit
      -- CP-element group 931: 	 branch_block_stmt_714/merge_stmt_2137_PhiAck/dummy
      -- 
    rr_5495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => type_cast_2141_inst_req_0); -- 
    cr_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => type_cast_2146_inst_req_1); -- 
    rr_5509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => type_cast_2146_inst_req_0); -- 
    cr_5500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => type_cast_2141_inst_req_1); -- 
    cr_5624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => ptr_deref_2190_store_0_req_1); -- 
    req_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => addr_of_2187_final_reg_req_1); -- 
    req_5559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => array_obj_ref_2186_index_offset_req_1); -- 
    cr_5528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(931), ack => type_cast_2180_inst_req_1); -- 
    zeropad3D_CP_2152_elements(931) <= OrReduce(zeropad3D_CP_2152_elements(253) & zeropad3D_CP_2152_elements(260) & zeropad3D_CP_2152_elements(263) & zeropad3D_CP_2152_elements(270));
    -- CP-element group 932:  merge  fork  transition  place  output  bypass 
    -- CP-element group 932: predecessors 
    -- CP-element group 932: 	284 
    -- CP-element group 932: 	304 
    -- CP-element group 932: successors 
    -- CP-element group 932: 	305 
    -- CP-element group 932: 	306 
    -- CP-element group 932:  members (13) 
      -- CP-element group 932: 	 branch_block_stmt_714/merge_stmt_2302__exit__
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320__entry__
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/$entry
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_sample_start_
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_update_start_
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Sample/$entry
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Sample/rr
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_714/assign_stmt_2307_to_assign_stmt_2320/type_cast_2306_Update/cr
      -- CP-element group 932: 	 branch_block_stmt_714/merge_stmt_2302_PhiReqMerge
      -- CP-element group 932: 	 branch_block_stmt_714/merge_stmt_2302_PhiAck/dummy
      -- CP-element group 932: 	 branch_block_stmt_714/merge_stmt_2302_PhiAck/$exit
      -- CP-element group 932: 	 branch_block_stmt_714/merge_stmt_2302_PhiAck/$entry
      -- 
    rr_5873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(932), ack => type_cast_2306_inst_req_0); -- 
    cr_5878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(932), ack => type_cast_2306_inst_req_1); -- 
    zeropad3D_CP_2152_elements(932) <= OrReduce(zeropad3D_CP_2152_elements(284) & zeropad3D_CP_2152_elements(304));
    -- CP-element group 933:  transition  output  delay-element  bypass 
    -- CP-element group 933: predecessors 
    -- CP-element group 933: 	326 
    -- CP-element group 933: successors 
    -- CP-element group 933: 	940 
    -- CP-element group 933:  members (4) 
      -- CP-element group 933: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_req
      -- CP-element group 933: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2427_konst_delay_trans
      -- CP-element group 933: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/$exit
      -- CP-element group 933: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2421/$exit
      -- 
    phi_stmt_2421_req_12445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2421_req_12445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(933), ack => phi_stmt_2421_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(933) is a control-delay.
    cp_element_933_delay: control_delay_element  generic map(name => " 933_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(326), ack => zeropad3D_CP_2152_elements(933), clk => clk, reset =>reset);
    -- CP-element group 934:  transition  input  bypass 
    -- CP-element group 934: predecessors 
    -- CP-element group 934: 	326 
    -- CP-element group 934: successors 
    -- CP-element group 934: 	936 
    -- CP-element group 934:  members (2) 
      -- CP-element group 934: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Sample/ra
      -- CP-element group 934: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Sample/$exit
      -- 
    ra_12462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 934_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2433_inst_ack_0, ack => zeropad3D_CP_2152_elements(934)); -- 
    -- CP-element group 935:  transition  input  bypass 
    -- CP-element group 935: predecessors 
    -- CP-element group 935: 	326 
    -- CP-element group 935: successors 
    -- CP-element group 935: 	936 
    -- CP-element group 935:  members (2) 
      -- CP-element group 935: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Update/ca
      -- CP-element group 935: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/Update/$exit
      -- 
    ca_12467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 935_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2433_inst_ack_1, ack => zeropad3D_CP_2152_elements(935)); -- 
    -- CP-element group 936:  join  transition  output  bypass 
    -- CP-element group 936: predecessors 
    -- CP-element group 936: 	934 
    -- CP-element group 936: 	935 
    -- CP-element group 936: successors 
    -- CP-element group 936: 	940 
    -- CP-element group 936:  members (5) 
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/$exit
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/$exit
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/SplitProtocol/$exit
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_req
      -- CP-element group 936: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2433/$exit
      -- 
    phi_stmt_2428_req_12468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2428_req_12468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(936), ack => phi_stmt_2428_req_1); -- 
    zeropad3D_cp_element_group_936: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_936"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(934) & zeropad3D_CP_2152_elements(935);
      gj_zeropad3D_cp_element_group_936 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(936), clk => clk, reset => reset); --
    end block;
    -- CP-element group 937:  transition  input  bypass 
    -- CP-element group 937: predecessors 
    -- CP-element group 937: 	326 
    -- CP-element group 937: successors 
    -- CP-element group 937: 	939 
    -- CP-element group 937:  members (2) 
      -- CP-element group 937: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Sample/ra
      -- CP-element group 937: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Sample/$exit
      -- 
    ra_12485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 937_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2439_inst_ack_0, ack => zeropad3D_CP_2152_elements(937)); -- 
    -- CP-element group 938:  transition  input  bypass 
    -- CP-element group 938: predecessors 
    -- CP-element group 938: 	326 
    -- CP-element group 938: successors 
    -- CP-element group 938: 	939 
    -- CP-element group 938:  members (2) 
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Update/ca
      -- CP-element group 938: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/Update/$exit
      -- 
    ca_12490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 938_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2439_inst_ack_1, ack => zeropad3D_CP_2152_elements(938)); -- 
    -- CP-element group 939:  join  transition  output  bypass 
    -- CP-element group 939: predecessors 
    -- CP-element group 939: 	937 
    -- CP-element group 939: 	938 
    -- CP-element group 939: successors 
    -- CP-element group 939: 	940 
    -- CP-element group 939:  members (5) 
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_req
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/SplitProtocol/$exit
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2439/$exit
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$exit
      -- CP-element group 939: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/phi_stmt_2434/$exit
      -- 
    phi_stmt_2434_req_12491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2434_req_12491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(939), ack => phi_stmt_2434_req_1); -- 
    zeropad3D_cp_element_group_939: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_939"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(937) & zeropad3D_CP_2152_elements(938);
      gj_zeropad3D_cp_element_group_939 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(939), clk => clk, reset => reset); --
    end block;
    -- CP-element group 940:  join  transition  bypass 
    -- CP-element group 940: predecessors 
    -- CP-element group 940: 	933 
    -- CP-element group 940: 	936 
    -- CP-element group 940: 	939 
    -- CP-element group 940: successors 
    -- CP-element group 940: 	951 
    -- CP-element group 940:  members (1) 
      -- CP-element group 940: 	 branch_block_stmt_714/ifx_xelse580_ifx_xend617_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_940: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_940"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(933) & zeropad3D_CP_2152_elements(936) & zeropad3D_CP_2152_elements(939);
      gj_zeropad3D_cp_element_group_940 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(940), clk => clk, reset => reset); --
    end block;
    -- CP-element group 941:  transition  input  bypass 
    -- CP-element group 941: predecessors 
    -- CP-element group 941: 	307 
    -- CP-element group 941: successors 
    -- CP-element group 941: 	943 
    -- CP-element group 941:  members (2) 
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Sample/ra
      -- CP-element group 941: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Sample/$exit
      -- 
    ra_12511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 941_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2424_inst_ack_0, ack => zeropad3D_CP_2152_elements(941)); -- 
    -- CP-element group 942:  transition  input  bypass 
    -- CP-element group 942: predecessors 
    -- CP-element group 942: 	307 
    -- CP-element group 942: successors 
    -- CP-element group 942: 	943 
    -- CP-element group 942:  members (2) 
      -- CP-element group 942: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Update/ca
      -- CP-element group 942: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/Update/$exit
      -- 
    ca_12516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 942_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2424_inst_ack_1, ack => zeropad3D_CP_2152_elements(942)); -- 
    -- CP-element group 943:  join  transition  output  bypass 
    -- CP-element group 943: predecessors 
    -- CP-element group 943: 	941 
    -- CP-element group 943: 	942 
    -- CP-element group 943: successors 
    -- CP-element group 943: 	950 
    -- CP-element group 943:  members (5) 
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/$exit
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_req
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/SplitProtocol/$exit
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/type_cast_2424/$exit
      -- CP-element group 943: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2421/phi_stmt_2421_sources/$exit
      -- 
    phi_stmt_2421_req_12517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2421_req_12517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(943), ack => phi_stmt_2421_req_0); -- 
    zeropad3D_cp_element_group_943: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_943"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(941) & zeropad3D_CP_2152_elements(942);
      gj_zeropad3D_cp_element_group_943 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(943), clk => clk, reset => reset); --
    end block;
    -- CP-element group 944:  transition  input  bypass 
    -- CP-element group 944: predecessors 
    -- CP-element group 944: 	307 
    -- CP-element group 944: successors 
    -- CP-element group 944: 	946 
    -- CP-element group 944:  members (2) 
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Sample/ra
      -- CP-element group 944: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Sample/$exit
      -- 
    ra_12534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 944_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_0, ack => zeropad3D_CP_2152_elements(944)); -- 
    -- CP-element group 945:  transition  input  bypass 
    -- CP-element group 945: predecessors 
    -- CP-element group 945: 	307 
    -- CP-element group 945: successors 
    -- CP-element group 945: 	946 
    -- CP-element group 945:  members (2) 
      -- CP-element group 945: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Update/ca
      -- CP-element group 945: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/Update/$exit
      -- 
    ca_12539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 945_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_1, ack => zeropad3D_CP_2152_elements(945)); -- 
    -- CP-element group 946:  join  transition  output  bypass 
    -- CP-element group 946: predecessors 
    -- CP-element group 946: 	944 
    -- CP-element group 946: 	945 
    -- CP-element group 946: successors 
    -- CP-element group 946: 	950 
    -- CP-element group 946:  members (5) 
      -- CP-element group 946: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/$exit
      -- CP-element group 946: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_req
      -- CP-element group 946: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/SplitProtocol/$exit
      -- CP-element group 946: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/type_cast_2431/$exit
      -- CP-element group 946: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2428/phi_stmt_2428_sources/$exit
      -- 
    phi_stmt_2428_req_12540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2428_req_12540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(946), ack => phi_stmt_2428_req_0); -- 
    zeropad3D_cp_element_group_946: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_946"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(944) & zeropad3D_CP_2152_elements(945);
      gj_zeropad3D_cp_element_group_946 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(946), clk => clk, reset => reset); --
    end block;
    -- CP-element group 947:  transition  input  bypass 
    -- CP-element group 947: predecessors 
    -- CP-element group 947: 	307 
    -- CP-element group 947: successors 
    -- CP-element group 947: 	949 
    -- CP-element group 947:  members (2) 
      -- CP-element group 947: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/ra
      -- CP-element group 947: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Sample/$exit
      -- 
    ra_12557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 947_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_0, ack => zeropad3D_CP_2152_elements(947)); -- 
    -- CP-element group 948:  transition  input  bypass 
    -- CP-element group 948: predecessors 
    -- CP-element group 948: 	307 
    -- CP-element group 948: successors 
    -- CP-element group 948: 	949 
    -- CP-element group 948:  members (2) 
      -- CP-element group 948: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/ca
      -- CP-element group 948: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/Update/$exit
      -- 
    ca_12562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 948_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_1, ack => zeropad3D_CP_2152_elements(948)); -- 
    -- CP-element group 949:  join  transition  output  bypass 
    -- CP-element group 949: predecessors 
    -- CP-element group 949: 	947 
    -- CP-element group 949: 	948 
    -- CP-element group 949: successors 
    -- CP-element group 949: 	950 
    -- CP-element group 949:  members (5) 
      -- CP-element group 949: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/SplitProtocol/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_req
      -- CP-element group 949: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/type_cast_2437/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/phi_stmt_2434_sources/$exit
      -- CP-element group 949: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/phi_stmt_2434/$exit
      -- 
    phi_stmt_2434_req_12563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2434_req_12563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(949), ack => phi_stmt_2434_req_0); -- 
    zeropad3D_cp_element_group_949: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_949"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(947) & zeropad3D_CP_2152_elements(948);
      gj_zeropad3D_cp_element_group_949 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(949), clk => clk, reset => reset); --
    end block;
    -- CP-element group 950:  join  transition  bypass 
    -- CP-element group 950: predecessors 
    -- CP-element group 950: 	943 
    -- CP-element group 950: 	946 
    -- CP-element group 950: 	949 
    -- CP-element group 950: successors 
    -- CP-element group 950: 	951 
    -- CP-element group 950:  members (1) 
      -- CP-element group 950: 	 branch_block_stmt_714/ifx_xthen575_ifx_xend617_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_950: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_950"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(943) & zeropad3D_CP_2152_elements(946) & zeropad3D_CP_2152_elements(949);
      gj_zeropad3D_cp_element_group_950 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(950), clk => clk, reset => reset); --
    end block;
    -- CP-element group 951:  merge  fork  transition  place  bypass 
    -- CP-element group 951: predecessors 
    -- CP-element group 951: 	940 
    -- CP-element group 951: 	950 
    -- CP-element group 951: successors 
    -- CP-element group 951: 	952 
    -- CP-element group 951: 	953 
    -- CP-element group 951: 	954 
    -- CP-element group 951:  members (2) 
      -- CP-element group 951: 	 branch_block_stmt_714/merge_stmt_2420_PhiAck/$entry
      -- CP-element group 951: 	 branch_block_stmt_714/merge_stmt_2420_PhiReqMerge
      -- 
    zeropad3D_CP_2152_elements(951) <= OrReduce(zeropad3D_CP_2152_elements(940) & zeropad3D_CP_2152_elements(950));
    -- CP-element group 952:  transition  input  bypass 
    -- CP-element group 952: predecessors 
    -- CP-element group 952: 	951 
    -- CP-element group 952: successors 
    -- CP-element group 952: 	955 
    -- CP-element group 952:  members (1) 
      -- CP-element group 952: 	 branch_block_stmt_714/merge_stmt_2420_PhiAck/phi_stmt_2421_ack
      -- 
    phi_stmt_2421_ack_12568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 952_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2421_ack_0, ack => zeropad3D_CP_2152_elements(952)); -- 
    -- CP-element group 953:  transition  input  bypass 
    -- CP-element group 953: predecessors 
    -- CP-element group 953: 	951 
    -- CP-element group 953: successors 
    -- CP-element group 953: 	955 
    -- CP-element group 953:  members (1) 
      -- CP-element group 953: 	 branch_block_stmt_714/merge_stmt_2420_PhiAck/phi_stmt_2428_ack
      -- 
    phi_stmt_2428_ack_12569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 953_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2428_ack_0, ack => zeropad3D_CP_2152_elements(953)); -- 
    -- CP-element group 954:  transition  input  bypass 
    -- CP-element group 954: predecessors 
    -- CP-element group 954: 	951 
    -- CP-element group 954: successors 
    -- CP-element group 954: 	955 
    -- CP-element group 954:  members (1) 
      -- CP-element group 954: 	 branch_block_stmt_714/merge_stmt_2420_PhiAck/phi_stmt_2434_ack
      -- 
    phi_stmt_2434_ack_12570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 954_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2434_ack_0, ack => zeropad3D_CP_2152_elements(954)); -- 
    -- CP-element group 955:  join  transition  bypass 
    -- CP-element group 955: predecessors 
    -- CP-element group 955: 	952 
    -- CP-element group 955: 	953 
    -- CP-element group 955: 	954 
    -- CP-element group 955: successors 
    -- CP-element group 955: 	3 
    -- CP-element group 955:  members (1) 
      -- CP-element group 955: 	 branch_block_stmt_714/merge_stmt_2420_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_955: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_955"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(952) & zeropad3D_CP_2152_elements(953) & zeropad3D_CP_2152_elements(954);
      gj_zeropad3D_cp_element_group_955 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(955), clk => clk, reset => reset); --
    end block;
    -- CP-element group 956:  transition  input  bypass 
    -- CP-element group 956: predecessors 
    -- CP-element group 956: 	4 
    -- CP-element group 956: successors 
    -- CP-element group 956: 	958 
    -- CP-element group 956:  members (2) 
      -- CP-element group 956: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Sample/$exit
      -- CP-element group 956: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Sample/ra
      -- 
    ra_12598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 956_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2596_inst_ack_0, ack => zeropad3D_CP_2152_elements(956)); -- 
    -- CP-element group 957:  transition  input  bypass 
    -- CP-element group 957: predecessors 
    -- CP-element group 957: 	4 
    -- CP-element group 957: successors 
    -- CP-element group 957: 	958 
    -- CP-element group 957:  members (2) 
      -- CP-element group 957: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Update/ca
      -- CP-element group 957: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/Update/$exit
      -- 
    ca_12603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 957_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2596_inst_ack_1, ack => zeropad3D_CP_2152_elements(957)); -- 
    -- CP-element group 958:  join  transition  output  bypass 
    -- CP-element group 958: predecessors 
    -- CP-element group 958: 	956 
    -- CP-element group 958: 	957 
    -- CP-element group 958: successors 
    -- CP-element group 958: 	965 
    -- CP-element group 958:  members (5) 
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/SplitProtocol/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2596/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/$exit
      -- CP-element group 958: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_req
      -- 
    phi_stmt_2590_req_12604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2590_req_12604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(958), ack => phi_stmt_2590_req_1); -- 
    zeropad3D_cp_element_group_958: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_958"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(956) & zeropad3D_CP_2152_elements(957);
      gj_zeropad3D_cp_element_group_958 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(958), clk => clk, reset => reset); --
    end block;
    -- CP-element group 959:  transition  input  bypass 
    -- CP-element group 959: predecessors 
    -- CP-element group 959: 	4 
    -- CP-element group 959: successors 
    -- CP-element group 959: 	961 
    -- CP-element group 959:  members (2) 
      -- CP-element group 959: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Sample/$exit
      -- CP-element group 959: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Sample/ra
      -- 
    ra_12621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 959_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2602_inst_ack_0, ack => zeropad3D_CP_2152_elements(959)); -- 
    -- CP-element group 960:  transition  input  bypass 
    -- CP-element group 960: predecessors 
    -- CP-element group 960: 	4 
    -- CP-element group 960: successors 
    -- CP-element group 960: 	961 
    -- CP-element group 960:  members (2) 
      -- CP-element group 960: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Update/ca
      -- CP-element group 960: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/Update/$exit
      -- 
    ca_12626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 960_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2602_inst_ack_1, ack => zeropad3D_CP_2152_elements(960)); -- 
    -- CP-element group 961:  join  transition  output  bypass 
    -- CP-element group 961: predecessors 
    -- CP-element group 961: 	959 
    -- CP-element group 961: 	960 
    -- CP-element group 961: successors 
    -- CP-element group 961: 	965 
    -- CP-element group 961:  members (5) 
      -- CP-element group 961: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_req
      -- CP-element group 961: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/SplitProtocol/$exit
      -- CP-element group 961: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2602/$exit
      -- CP-element group 961: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/$exit
      -- CP-element group 961: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2597/$exit
      -- 
    phi_stmt_2597_req_12627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2597_req_12627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(961), ack => phi_stmt_2597_req_1); -- 
    zeropad3D_cp_element_group_961: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_961"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(959) & zeropad3D_CP_2152_elements(960);
      gj_zeropad3D_cp_element_group_961 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(961), clk => clk, reset => reset); --
    end block;
    -- CP-element group 962:  transition  input  bypass 
    -- CP-element group 962: predecessors 
    -- CP-element group 962: 	4 
    -- CP-element group 962: successors 
    -- CP-element group 962: 	964 
    -- CP-element group 962:  members (2) 
      -- CP-element group 962: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Sample/$exit
      -- CP-element group 962: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Sample/ra
      -- 
    ra_12644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 962_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2608_inst_ack_0, ack => zeropad3D_CP_2152_elements(962)); -- 
    -- CP-element group 963:  transition  input  bypass 
    -- CP-element group 963: predecessors 
    -- CP-element group 963: 	4 
    -- CP-element group 963: successors 
    -- CP-element group 963: 	964 
    -- CP-element group 963:  members (2) 
      -- CP-element group 963: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Update/$exit
      -- CP-element group 963: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/Update/ca
      -- 
    ca_12649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 963_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2608_inst_ack_1, ack => zeropad3D_CP_2152_elements(963)); -- 
    -- CP-element group 964:  join  transition  output  bypass 
    -- CP-element group 964: predecessors 
    -- CP-element group 964: 	962 
    -- CP-element group 964: 	963 
    -- CP-element group 964: successors 
    -- CP-element group 964: 	965 
    -- CP-element group 964:  members (5) 
      -- CP-element group 964: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/$exit
      -- CP-element group 964: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$exit
      -- CP-element group 964: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/$exit
      -- CP-element group 964: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2608/SplitProtocol/$exit
      -- CP-element group 964: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_req
      -- 
    phi_stmt_2603_req_12650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2603_req_12650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(964), ack => phi_stmt_2603_req_1); -- 
    zeropad3D_cp_element_group_964: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_964"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(962) & zeropad3D_CP_2152_elements(963);
      gj_zeropad3D_cp_element_group_964 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(964), clk => clk, reset => reset); --
    end block;
    -- CP-element group 965:  join  transition  bypass 
    -- CP-element group 965: predecessors 
    -- CP-element group 965: 	958 
    -- CP-element group 965: 	961 
    -- CP-element group 965: 	964 
    -- CP-element group 965: successors 
    -- CP-element group 965: 	974 
    -- CP-element group 965:  members (1) 
      -- CP-element group 965: 	 branch_block_stmt_714/ifx_xend837_whilex_xbody682_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_965: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_965"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(958) & zeropad3D_CP_2152_elements(961) & zeropad3D_CP_2152_elements(964);
      gj_zeropad3D_cp_element_group_965 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(965), clk => clk, reset => reset); --
    end block;
    -- CP-element group 966:  transition  output  delay-element  bypass 
    -- CP-element group 966: predecessors 
    -- CP-element group 966: 	349 
    -- CP-element group 966: successors 
    -- CP-element group 966: 	973 
    -- CP-element group 966:  members (4) 
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2590/$exit
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/$exit
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_sources/type_cast_2594_konst_delay_trans
      -- CP-element group 966: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2590/phi_stmt_2590_req
      -- 
    phi_stmt_2590_req_12661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2590_req_12661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(966), ack => phi_stmt_2590_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(966) is a control-delay.
    cp_element_966_delay: control_delay_element  generic map(name => " 966_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(349), ack => zeropad3D_CP_2152_elements(966), clk => clk, reset =>reset);
    -- CP-element group 967:  transition  input  bypass 
    -- CP-element group 967: predecessors 
    -- CP-element group 967: 	349 
    -- CP-element group 967: successors 
    -- CP-element group 967: 	969 
    -- CP-element group 967:  members (2) 
      -- CP-element group 967: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Sample/$exit
      -- CP-element group 967: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Sample/ra
      -- 
    ra_12678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 967_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2600_inst_ack_0, ack => zeropad3D_CP_2152_elements(967)); -- 
    -- CP-element group 968:  transition  input  bypass 
    -- CP-element group 968: predecessors 
    -- CP-element group 968: 	349 
    -- CP-element group 968: successors 
    -- CP-element group 968: 	969 
    -- CP-element group 968:  members (2) 
      -- CP-element group 968: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Update/$exit
      -- CP-element group 968: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/Update/ca
      -- 
    ca_12683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 968_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2600_inst_ack_1, ack => zeropad3D_CP_2152_elements(968)); -- 
    -- CP-element group 969:  join  transition  output  bypass 
    -- CP-element group 969: predecessors 
    -- CP-element group 969: 	967 
    -- CP-element group 969: 	968 
    -- CP-element group 969: successors 
    -- CP-element group 969: 	973 
    -- CP-element group 969:  members (5) 
      -- CP-element group 969: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/$exit
      -- CP-element group 969: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/$exit
      -- CP-element group 969: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/$exit
      -- CP-element group 969: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_sources/type_cast_2600/SplitProtocol/$exit
      -- CP-element group 969: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2597/phi_stmt_2597_req
      -- 
    phi_stmt_2597_req_12684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2597_req_12684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(969), ack => phi_stmt_2597_req_0); -- 
    zeropad3D_cp_element_group_969: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_969"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(967) & zeropad3D_CP_2152_elements(968);
      gj_zeropad3D_cp_element_group_969 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(969), clk => clk, reset => reset); --
    end block;
    -- CP-element group 970:  transition  input  bypass 
    -- CP-element group 970: predecessors 
    -- CP-element group 970: 	349 
    -- CP-element group 970: successors 
    -- CP-element group 970: 	972 
    -- CP-element group 970:  members (2) 
      -- CP-element group 970: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Sample/$exit
      -- CP-element group 970: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Sample/ra
      -- 
    ra_12701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 970_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_0, ack => zeropad3D_CP_2152_elements(970)); -- 
    -- CP-element group 971:  transition  input  bypass 
    -- CP-element group 971: predecessors 
    -- CP-element group 971: 	349 
    -- CP-element group 971: successors 
    -- CP-element group 971: 	972 
    -- CP-element group 971:  members (2) 
      -- CP-element group 971: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Update/$exit
      -- CP-element group 971: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/Update/ca
      -- 
    ca_12706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 971_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_1, ack => zeropad3D_CP_2152_elements(971)); -- 
    -- CP-element group 972:  join  transition  output  bypass 
    -- CP-element group 972: predecessors 
    -- CP-element group 972: 	970 
    -- CP-element group 972: 	971 
    -- CP-element group 972: successors 
    -- CP-element group 972: 	973 
    -- CP-element group 972:  members (5) 
      -- CP-element group 972: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/$exit
      -- CP-element group 972: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$exit
      -- CP-element group 972: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/$exit
      -- CP-element group 972: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2606/SplitProtocol/$exit
      -- CP-element group 972: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/phi_stmt_2603/phi_stmt_2603_req
      -- 
    phi_stmt_2603_req_12707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2603_req_12707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(972), ack => phi_stmt_2603_req_0); -- 
    zeropad3D_cp_element_group_972: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_972"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(970) & zeropad3D_CP_2152_elements(971);
      gj_zeropad3D_cp_element_group_972 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(972), clk => clk, reset => reset); --
    end block;
    -- CP-element group 973:  join  transition  bypass 
    -- CP-element group 973: predecessors 
    -- CP-element group 973: 	966 
    -- CP-element group 973: 	969 
    -- CP-element group 973: 	972 
    -- CP-element group 973: successors 
    -- CP-element group 973: 	974 
    -- CP-element group 973:  members (1) 
      -- CP-element group 973: 	 branch_block_stmt_714/whilex_xend618_whilex_xbody682_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_973: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_973"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(966) & zeropad3D_CP_2152_elements(969) & zeropad3D_CP_2152_elements(972);
      gj_zeropad3D_cp_element_group_973 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(973), clk => clk, reset => reset); --
    end block;
    -- CP-element group 974:  merge  fork  transition  place  bypass 
    -- CP-element group 974: predecessors 
    -- CP-element group 974: 	965 
    -- CP-element group 974: 	973 
    -- CP-element group 974: successors 
    -- CP-element group 974: 	975 
    -- CP-element group 974: 	976 
    -- CP-element group 974: 	977 
    -- CP-element group 974:  members (2) 
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2589_PhiReqMerge
      -- CP-element group 974: 	 branch_block_stmt_714/merge_stmt_2589_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(974) <= OrReduce(zeropad3D_CP_2152_elements(965) & zeropad3D_CP_2152_elements(973));
    -- CP-element group 975:  transition  input  bypass 
    -- CP-element group 975: predecessors 
    -- CP-element group 975: 	974 
    -- CP-element group 975: successors 
    -- CP-element group 975: 	978 
    -- CP-element group 975:  members (1) 
      -- CP-element group 975: 	 branch_block_stmt_714/merge_stmt_2589_PhiAck/phi_stmt_2590_ack
      -- 
    phi_stmt_2590_ack_12712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 975_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2590_ack_0, ack => zeropad3D_CP_2152_elements(975)); -- 
    -- CP-element group 976:  transition  input  bypass 
    -- CP-element group 976: predecessors 
    -- CP-element group 976: 	974 
    -- CP-element group 976: successors 
    -- CP-element group 976: 	978 
    -- CP-element group 976:  members (1) 
      -- CP-element group 976: 	 branch_block_stmt_714/merge_stmt_2589_PhiAck/phi_stmt_2597_ack
      -- 
    phi_stmt_2597_ack_12713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 976_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2597_ack_0, ack => zeropad3D_CP_2152_elements(976)); -- 
    -- CP-element group 977:  transition  input  bypass 
    -- CP-element group 977: predecessors 
    -- CP-element group 977: 	974 
    -- CP-element group 977: successors 
    -- CP-element group 977: 	978 
    -- CP-element group 977:  members (1) 
      -- CP-element group 977: 	 branch_block_stmt_714/merge_stmt_2589_PhiAck/phi_stmt_2603_ack
      -- 
    phi_stmt_2603_ack_12714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 977_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2603_ack_0, ack => zeropad3D_CP_2152_elements(977)); -- 
    -- CP-element group 978:  join  fork  transition  place  output  bypass 
    -- CP-element group 978: predecessors 
    -- CP-element group 978: 	975 
    -- CP-element group 978: 	976 
    -- CP-element group 978: 	977 
    -- CP-element group 978: successors 
    -- CP-element group 978: 	350 
    -- CP-element group 978: 	351 
    -- CP-element group 978:  members (10) 
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621__entry__
      -- CP-element group 978: 	 branch_block_stmt_714/merge_stmt_2589__exit__
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/$entry
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_sample_start_
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_update_start_
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Sample/$entry
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Sample/rr
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Update/$entry
      -- CP-element group 978: 	 branch_block_stmt_714/assign_stmt_2614_to_assign_stmt_2621/type_cast_2613_Update/cr
      -- CP-element group 978: 	 branch_block_stmt_714/merge_stmt_2589_PhiAck/$exit
      -- 
    rr_6375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(978), ack => type_cast_2613_inst_req_0); -- 
    cr_6380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(978), ack => type_cast_2613_inst_req_1); -- 
    zeropad3D_cp_element_group_978: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_978"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(975) & zeropad3D_CP_2152_elements(976) & zeropad3D_CP_2152_elements(977);
      gj_zeropad3D_cp_element_group_978 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(978), clk => clk, reset => reset); --
    end block;
    -- CP-element group 979:  merge  fork  transition  place  output  bypass 
    -- CP-element group 979: predecessors 
    -- CP-element group 979: 	352 
    -- CP-element group 979: 	359 
    -- CP-element group 979: 	362 
    -- CP-element group 979: 	369 
    -- CP-element group 979: successors 
    -- CP-element group 979: 	370 
    -- CP-element group 979: 	371 
    -- CP-element group 979: 	372 
    -- CP-element group 979: 	373 
    -- CP-element group 979: 	376 
    -- CP-element group 979: 	378 
    -- CP-element group 979: 	380 
    -- CP-element group 979: 	382 
    -- CP-element group 979:  members (33) 
      -- CP-element group 979: 	 branch_block_stmt_714/merge_stmt_2705__exit__
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761__entry__
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Update/req
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_Update/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_update_start_
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/array_obj_ref_2754_final_index_sum_regn_update_start
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/word_access_complete/word_0/cr
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/word_access_complete/word_0/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/word_access_complete/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_complete/req
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/ptr_deref_2758_Update/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_complete/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_sample_start_
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_update_start_
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Sample/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Sample/rr
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Update/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2709_Update/cr
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_sample_start_
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_update_start_
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Sample/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Sample/rr
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Update/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2714_Update/cr
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_update_start_
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Update/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/type_cast_2748_Update/cr
      -- CP-element group 979: 	 branch_block_stmt_714/assign_stmt_2710_to_assign_stmt_2761/addr_of_2755_update_start_
      -- CP-element group 979: 	 branch_block_stmt_714/merge_stmt_2705_PhiReqMerge
      -- CP-element group 979: 	 branch_block_stmt_714/merge_stmt_2705_PhiAck/$entry
      -- CP-element group 979: 	 branch_block_stmt_714/merge_stmt_2705_PhiAck/$exit
      -- CP-element group 979: 	 branch_block_stmt_714/merge_stmt_2705_PhiAck/dummy
      -- 
    req_6649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => array_obj_ref_2754_index_offset_req_1); -- 
    cr_6714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => ptr_deref_2758_store_0_req_1); -- 
    req_6664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => addr_of_2755_final_reg_req_1); -- 
    rr_6585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => type_cast_2709_inst_req_0); -- 
    cr_6590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => type_cast_2709_inst_req_1); -- 
    rr_6599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => type_cast_2714_inst_req_0); -- 
    cr_6604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => type_cast_2714_inst_req_1); -- 
    cr_6618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(979), ack => type_cast_2748_inst_req_1); -- 
    zeropad3D_CP_2152_elements(979) <= OrReduce(zeropad3D_CP_2152_elements(352) & zeropad3D_CP_2152_elements(359) & zeropad3D_CP_2152_elements(362) & zeropad3D_CP_2152_elements(369));
    -- CP-element group 980:  merge  fork  transition  place  output  bypass 
    -- CP-element group 980: predecessors 
    -- CP-element group 980: 	383 
    -- CP-element group 980: 	403 
    -- CP-element group 980: successors 
    -- CP-element group 980: 	404 
    -- CP-element group 980: 	405 
    -- CP-element group 980:  members (13) 
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888__entry__
      -- CP-element group 980: 	 branch_block_stmt_714/merge_stmt_2870__exit__
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/$entry
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_sample_start_
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_update_start_
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Sample/$entry
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Sample/rr
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Update/$entry
      -- CP-element group 980: 	 branch_block_stmt_714/assign_stmt_2875_to_assign_stmt_2888/type_cast_2874_Update/cr
      -- CP-element group 980: 	 branch_block_stmt_714/merge_stmt_2870_PhiReqMerge
      -- CP-element group 980: 	 branch_block_stmt_714/merge_stmt_2870_PhiAck/$entry
      -- CP-element group 980: 	 branch_block_stmt_714/merge_stmt_2870_PhiAck/$exit
      -- CP-element group 980: 	 branch_block_stmt_714/merge_stmt_2870_PhiAck/dummy
      -- 
    rr_6963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(980), ack => type_cast_2874_inst_req_0); -- 
    cr_6968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(980), ack => type_cast_2874_inst_req_1); -- 
    zeropad3D_CP_2152_elements(980) <= OrReduce(zeropad3D_CP_2152_elements(383) & zeropad3D_CP_2152_elements(403));
    -- CP-element group 981:  transition  output  delay-element  bypass 
    -- CP-element group 981: predecessors 
    -- CP-element group 981: 	425 
    -- CP-element group 981: successors 
    -- CP-element group 981: 	988 
    -- CP-element group 981:  members (4) 
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2982/$exit
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/$exit
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2988_konst_delay_trans
      -- CP-element group 981: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_req
      -- 
    phi_stmt_2982_req_12825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2982_req_12825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(981), ack => phi_stmt_2982_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(981) is a control-delay.
    cp_element_981_delay: control_delay_element  generic map(name => " 981_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(425), ack => zeropad3D_CP_2152_elements(981), clk => clk, reset =>reset);
    -- CP-element group 982:  transition  input  bypass 
    -- CP-element group 982: predecessors 
    -- CP-element group 982: 	425 
    -- CP-element group 982: successors 
    -- CP-element group 982: 	984 
    -- CP-element group 982:  members (2) 
      -- CP-element group 982: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Sample/$exit
      -- CP-element group 982: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Sample/ra
      -- 
    ra_12842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 982_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2994_inst_ack_0, ack => zeropad3D_CP_2152_elements(982)); -- 
    -- CP-element group 983:  transition  input  bypass 
    -- CP-element group 983: predecessors 
    -- CP-element group 983: 	425 
    -- CP-element group 983: successors 
    -- CP-element group 983: 	984 
    -- CP-element group 983:  members (2) 
      -- CP-element group 983: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Update/$exit
      -- CP-element group 983: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/Update/ca
      -- 
    ca_12847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 983_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2994_inst_ack_1, ack => zeropad3D_CP_2152_elements(983)); -- 
    -- CP-element group 984:  join  transition  output  bypass 
    -- CP-element group 984: predecessors 
    -- CP-element group 984: 	982 
    -- CP-element group 984: 	983 
    -- CP-element group 984: successors 
    -- CP-element group 984: 	988 
    -- CP-element group 984:  members (5) 
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/$exit
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/$exit
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/$exit
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2994/SplitProtocol/$exit
      -- CP-element group 984: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_req
      -- 
    phi_stmt_2989_req_12848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2989_req_12848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(984), ack => phi_stmt_2989_req_1); -- 
    zeropad3D_cp_element_group_984: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_984"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(982) & zeropad3D_CP_2152_elements(983);
      gj_zeropad3D_cp_element_group_984 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(984), clk => clk, reset => reset); --
    end block;
    -- CP-element group 985:  transition  input  bypass 
    -- CP-element group 985: predecessors 
    -- CP-element group 985: 	425 
    -- CP-element group 985: successors 
    -- CP-element group 985: 	987 
    -- CP-element group 985:  members (2) 
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Sample/$exit
      -- CP-element group 985: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Sample/ra
      -- 
    ra_12865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 985_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3000_inst_ack_0, ack => zeropad3D_CP_2152_elements(985)); -- 
    -- CP-element group 986:  transition  input  bypass 
    -- CP-element group 986: predecessors 
    -- CP-element group 986: 	425 
    -- CP-element group 986: successors 
    -- CP-element group 986: 	987 
    -- CP-element group 986:  members (2) 
      -- CP-element group 986: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Update/$exit
      -- CP-element group 986: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/Update/ca
      -- 
    ca_12870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 986_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3000_inst_ack_1, ack => zeropad3D_CP_2152_elements(986)); -- 
    -- CP-element group 987:  join  transition  output  bypass 
    -- CP-element group 987: predecessors 
    -- CP-element group 987: 	985 
    -- CP-element group 987: 	986 
    -- CP-element group 987: successors 
    -- CP-element group 987: 	988 
    -- CP-element group 987:  members (5) 
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/$exit
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/$exit
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/$exit
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_3000/SplitProtocol/$exit
      -- CP-element group 987: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_req
      -- 
    phi_stmt_2995_req_12871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2995_req_12871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(987), ack => phi_stmt_2995_req_1); -- 
    zeropad3D_cp_element_group_987: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_987"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(985) & zeropad3D_CP_2152_elements(986);
      gj_zeropad3D_cp_element_group_987 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(987), clk => clk, reset => reset); --
    end block;
    -- CP-element group 988:  join  transition  bypass 
    -- CP-element group 988: predecessors 
    -- CP-element group 988: 	981 
    -- CP-element group 988: 	984 
    -- CP-element group 988: 	987 
    -- CP-element group 988: successors 
    -- CP-element group 988: 	999 
    -- CP-element group 988:  members (1) 
      -- CP-element group 988: 	 branch_block_stmt_714/ifx_xelse801_ifx_xend837_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_988: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_988"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(981) & zeropad3D_CP_2152_elements(984) & zeropad3D_CP_2152_elements(987);
      gj_zeropad3D_cp_element_group_988 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(988), clk => clk, reset => reset); --
    end block;
    -- CP-element group 989:  transition  input  bypass 
    -- CP-element group 989: predecessors 
    -- CP-element group 989: 	406 
    -- CP-element group 989: successors 
    -- CP-element group 989: 	991 
    -- CP-element group 989:  members (2) 
      -- CP-element group 989: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Sample/$exit
      -- CP-element group 989: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Sample/ra
      -- 
    ra_12891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 989_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2985_inst_ack_0, ack => zeropad3D_CP_2152_elements(989)); -- 
    -- CP-element group 990:  transition  input  bypass 
    -- CP-element group 990: predecessors 
    -- CP-element group 990: 	406 
    -- CP-element group 990: successors 
    -- CP-element group 990: 	991 
    -- CP-element group 990:  members (2) 
      -- CP-element group 990: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Update/$exit
      -- CP-element group 990: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/Update/ca
      -- 
    ca_12896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 990_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2985_inst_ack_1, ack => zeropad3D_CP_2152_elements(990)); -- 
    -- CP-element group 991:  join  transition  output  bypass 
    -- CP-element group 991: predecessors 
    -- CP-element group 991: 	989 
    -- CP-element group 991: 	990 
    -- CP-element group 991: successors 
    -- CP-element group 991: 	998 
    -- CP-element group 991:  members (5) 
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_sources/type_cast_2985/SplitProtocol/$exit
      -- CP-element group 991: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2982/phi_stmt_2982_req
      -- 
    phi_stmt_2982_req_12897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2982_req_12897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(991), ack => phi_stmt_2982_req_0); -- 
    zeropad3D_cp_element_group_991: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_991"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(989) & zeropad3D_CP_2152_elements(990);
      gj_zeropad3D_cp_element_group_991 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(991), clk => clk, reset => reset); --
    end block;
    -- CP-element group 992:  transition  input  bypass 
    -- CP-element group 992: predecessors 
    -- CP-element group 992: 	406 
    -- CP-element group 992: successors 
    -- CP-element group 992: 	994 
    -- CP-element group 992:  members (2) 
      -- CP-element group 992: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Sample/$exit
      -- CP-element group 992: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Sample/ra
      -- 
    ra_12914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 992_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2992_inst_ack_0, ack => zeropad3D_CP_2152_elements(992)); -- 
    -- CP-element group 993:  transition  input  bypass 
    -- CP-element group 993: predecessors 
    -- CP-element group 993: 	406 
    -- CP-element group 993: successors 
    -- CP-element group 993: 	994 
    -- CP-element group 993:  members (2) 
      -- CP-element group 993: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Update/$exit
      -- CP-element group 993: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/Update/ca
      -- 
    ca_12919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 993_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2992_inst_ack_1, ack => zeropad3D_CP_2152_elements(993)); -- 
    -- CP-element group 994:  join  transition  output  bypass 
    -- CP-element group 994: predecessors 
    -- CP-element group 994: 	992 
    -- CP-element group 994: 	993 
    -- CP-element group 994: successors 
    -- CP-element group 994: 	998 
    -- CP-element group 994:  members (5) 
      -- CP-element group 994: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/$exit
      -- CP-element group 994: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/$exit
      -- CP-element group 994: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/$exit
      -- CP-element group 994: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_sources/type_cast_2992/SplitProtocol/$exit
      -- CP-element group 994: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2989/phi_stmt_2989_req
      -- 
    phi_stmt_2989_req_12920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2989_req_12920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(994), ack => phi_stmt_2989_req_0); -- 
    zeropad3D_cp_element_group_994: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_994"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(992) & zeropad3D_CP_2152_elements(993);
      gj_zeropad3D_cp_element_group_994 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(994), clk => clk, reset => reset); --
    end block;
    -- CP-element group 995:  transition  input  bypass 
    -- CP-element group 995: predecessors 
    -- CP-element group 995: 	406 
    -- CP-element group 995: successors 
    -- CP-element group 995: 	997 
    -- CP-element group 995:  members (2) 
      -- CP-element group 995: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Sample/$exit
      -- CP-element group 995: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Sample/ra
      -- 
    ra_12937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 995_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2998_inst_ack_0, ack => zeropad3D_CP_2152_elements(995)); -- 
    -- CP-element group 996:  transition  input  bypass 
    -- CP-element group 996: predecessors 
    -- CP-element group 996: 	406 
    -- CP-element group 996: successors 
    -- CP-element group 996: 	997 
    -- CP-element group 996:  members (2) 
      -- CP-element group 996: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Update/$exit
      -- CP-element group 996: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/Update/ca
      -- 
    ca_12942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 996_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2998_inst_ack_1, ack => zeropad3D_CP_2152_elements(996)); -- 
    -- CP-element group 997:  join  transition  output  bypass 
    -- CP-element group 997: predecessors 
    -- CP-element group 997: 	995 
    -- CP-element group 997: 	996 
    -- CP-element group 997: successors 
    -- CP-element group 997: 	998 
    -- CP-element group 997:  members (5) 
      -- CP-element group 997: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/$exit
      -- CP-element group 997: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/$exit
      -- CP-element group 997: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/$exit
      -- CP-element group 997: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_sources/type_cast_2998/SplitProtocol/$exit
      -- CP-element group 997: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/phi_stmt_2995/phi_stmt_2995_req
      -- 
    phi_stmt_2995_req_12943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2995_req_12943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(997), ack => phi_stmt_2995_req_0); -- 
    zeropad3D_cp_element_group_997: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_997"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(995) & zeropad3D_CP_2152_elements(996);
      gj_zeropad3D_cp_element_group_997 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(997), clk => clk, reset => reset); --
    end block;
    -- CP-element group 998:  join  transition  bypass 
    -- CP-element group 998: predecessors 
    -- CP-element group 998: 	991 
    -- CP-element group 998: 	994 
    -- CP-element group 998: 	997 
    -- CP-element group 998: successors 
    -- CP-element group 998: 	999 
    -- CP-element group 998:  members (1) 
      -- CP-element group 998: 	 branch_block_stmt_714/ifx_xthen796_ifx_xend837_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_998: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_998"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(991) & zeropad3D_CP_2152_elements(994) & zeropad3D_CP_2152_elements(997);
      gj_zeropad3D_cp_element_group_998 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(998), clk => clk, reset => reset); --
    end block;
    -- CP-element group 999:  merge  fork  transition  place  bypass 
    -- CP-element group 999: predecessors 
    -- CP-element group 999: 	988 
    -- CP-element group 999: 	998 
    -- CP-element group 999: successors 
    -- CP-element group 999: 	1000 
    -- CP-element group 999: 	1001 
    -- CP-element group 999: 	1002 
    -- CP-element group 999:  members (2) 
      -- CP-element group 999: 	 branch_block_stmt_714/merge_stmt_2981_PhiReqMerge
      -- CP-element group 999: 	 branch_block_stmt_714/merge_stmt_2981_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(999) <= OrReduce(zeropad3D_CP_2152_elements(988) & zeropad3D_CP_2152_elements(998));
    -- CP-element group 1000:  transition  input  bypass 
    -- CP-element group 1000: predecessors 
    -- CP-element group 1000: 	999 
    -- CP-element group 1000: successors 
    -- CP-element group 1000: 	1003 
    -- CP-element group 1000:  members (1) 
      -- CP-element group 1000: 	 branch_block_stmt_714/merge_stmt_2981_PhiAck/phi_stmt_2982_ack
      -- 
    phi_stmt_2982_ack_12948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1000_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2982_ack_0, ack => zeropad3D_CP_2152_elements(1000)); -- 
    -- CP-element group 1001:  transition  input  bypass 
    -- CP-element group 1001: predecessors 
    -- CP-element group 1001: 	999 
    -- CP-element group 1001: successors 
    -- CP-element group 1001: 	1003 
    -- CP-element group 1001:  members (1) 
      -- CP-element group 1001: 	 branch_block_stmt_714/merge_stmt_2981_PhiAck/phi_stmt_2989_ack
      -- 
    phi_stmt_2989_ack_12949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1001_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2989_ack_0, ack => zeropad3D_CP_2152_elements(1001)); -- 
    -- CP-element group 1002:  transition  input  bypass 
    -- CP-element group 1002: predecessors 
    -- CP-element group 1002: 	999 
    -- CP-element group 1002: successors 
    -- CP-element group 1002: 	1003 
    -- CP-element group 1002:  members (1) 
      -- CP-element group 1002: 	 branch_block_stmt_714/merge_stmt_2981_PhiAck/phi_stmt_2995_ack
      -- 
    phi_stmt_2995_ack_12950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1002_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2995_ack_0, ack => zeropad3D_CP_2152_elements(1002)); -- 
    -- CP-element group 1003:  join  transition  bypass 
    -- CP-element group 1003: predecessors 
    -- CP-element group 1003: 	1000 
    -- CP-element group 1003: 	1001 
    -- CP-element group 1003: 	1002 
    -- CP-element group 1003: successors 
    -- CP-element group 1003: 	4 
    -- CP-element group 1003:  members (1) 
      -- CP-element group 1003: 	 branch_block_stmt_714/merge_stmt_2981_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1003: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1003"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1000) & zeropad3D_CP_2152_elements(1001) & zeropad3D_CP_2152_elements(1002);
      gj_zeropad3D_cp_element_group_1003 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1003), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1004:  transition  input  bypass 
    -- CP-element group 1004: predecessors 
    -- CP-element group 1004: 	5 
    -- CP-element group 1004: successors 
    -- CP-element group 1004: 	1006 
    -- CP-element group 1004:  members (2) 
      -- CP-element group 1004: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Sample/$exit
      -- CP-element group 1004: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Sample/ra
      -- 
    ra_12978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1004_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3157_inst_ack_0, ack => zeropad3D_CP_2152_elements(1004)); -- 
    -- CP-element group 1005:  transition  input  bypass 
    -- CP-element group 1005: predecessors 
    -- CP-element group 1005: 	5 
    -- CP-element group 1005: successors 
    -- CP-element group 1005: 	1006 
    -- CP-element group 1005:  members (2) 
      -- CP-element group 1005: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Update/$exit
      -- CP-element group 1005: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/Update/ca
      -- 
    ca_12983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1005_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3157_inst_ack_1, ack => zeropad3D_CP_2152_elements(1005)); -- 
    -- CP-element group 1006:  join  transition  output  bypass 
    -- CP-element group 1006: predecessors 
    -- CP-element group 1006: 	1004 
    -- CP-element group 1006: 	1005 
    -- CP-element group 1006: successors 
    -- CP-element group 1006: 	1013 
    -- CP-element group 1006:  members (5) 
      -- CP-element group 1006: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/$exit
      -- CP-element group 1006: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/$exit
      -- CP-element group 1006: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/$exit
      -- CP-element group 1006: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3157/SplitProtocol/$exit
      -- CP-element group 1006: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_req
      -- 
    phi_stmt_3154_req_12984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3154_req_12984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1006), ack => phi_stmt_3154_req_0); -- 
    zeropad3D_cp_element_group_1006: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1006"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1004) & zeropad3D_CP_2152_elements(1005);
      gj_zeropad3D_cp_element_group_1006 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1006), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1007:  transition  input  bypass 
    -- CP-element group 1007: predecessors 
    -- CP-element group 1007: 	5 
    -- CP-element group 1007: successors 
    -- CP-element group 1007: 	1009 
    -- CP-element group 1007:  members (2) 
      -- CP-element group 1007: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Sample/$exit
      -- CP-element group 1007: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Sample/ra
      -- 
    ra_13001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1007_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3153_inst_ack_0, ack => zeropad3D_CP_2152_elements(1007)); -- 
    -- CP-element group 1008:  transition  input  bypass 
    -- CP-element group 1008: predecessors 
    -- CP-element group 1008: 	5 
    -- CP-element group 1008: successors 
    -- CP-element group 1008: 	1009 
    -- CP-element group 1008:  members (2) 
      -- CP-element group 1008: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Update/$exit
      -- CP-element group 1008: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/Update/ca
      -- 
    ca_13006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1008_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3153_inst_ack_1, ack => zeropad3D_CP_2152_elements(1008)); -- 
    -- CP-element group 1009:  join  transition  output  bypass 
    -- CP-element group 1009: predecessors 
    -- CP-element group 1009: 	1007 
    -- CP-element group 1009: 	1008 
    -- CP-element group 1009: successors 
    -- CP-element group 1009: 	1013 
    -- CP-element group 1009:  members (5) 
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/$exit
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/$exit
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/$exit
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3153/SplitProtocol/$exit
      -- CP-element group 1009: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_req
      -- 
    phi_stmt_3148_req_13007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3148_req_13007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1009), ack => phi_stmt_3148_req_1); -- 
    zeropad3D_cp_element_group_1009: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1009"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1007) & zeropad3D_CP_2152_elements(1008);
      gj_zeropad3D_cp_element_group_1009 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1009), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1010:  transition  input  bypass 
    -- CP-element group 1010: predecessors 
    -- CP-element group 1010: 	5 
    -- CP-element group 1010: successors 
    -- CP-element group 1010: 	1012 
    -- CP-element group 1010:  members (2) 
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Sample/$exit
      -- CP-element group 1010: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Sample/ra
      -- 
    ra_13024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1010_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3144_inst_ack_0, ack => zeropad3D_CP_2152_elements(1010)); -- 
    -- CP-element group 1011:  transition  input  bypass 
    -- CP-element group 1011: predecessors 
    -- CP-element group 1011: 	5 
    -- CP-element group 1011: successors 
    -- CP-element group 1011: 	1012 
    -- CP-element group 1011:  members (2) 
      -- CP-element group 1011: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Update/$exit
      -- CP-element group 1011: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/Update/ca
      -- 
    ca_13029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1011_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3144_inst_ack_1, ack => zeropad3D_CP_2152_elements(1011)); -- 
    -- CP-element group 1012:  join  transition  output  bypass 
    -- CP-element group 1012: predecessors 
    -- CP-element group 1012: 	1010 
    -- CP-element group 1012: 	1011 
    -- CP-element group 1012: successors 
    -- CP-element group 1012: 	1013 
    -- CP-element group 1012:  members (5) 
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/$exit
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/$exit
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/$exit
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3144/SplitProtocol/$exit
      -- CP-element group 1012: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_req
      -- 
    phi_stmt_3141_req_13030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3141_req_13030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1012), ack => phi_stmt_3141_req_0); -- 
    zeropad3D_cp_element_group_1012: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1012"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1010) & zeropad3D_CP_2152_elements(1011);
      gj_zeropad3D_cp_element_group_1012 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1012), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1013:  join  transition  bypass 
    -- CP-element group 1013: predecessors 
    -- CP-element group 1013: 	1006 
    -- CP-element group 1013: 	1009 
    -- CP-element group 1013: 	1012 
    -- CP-element group 1013: successors 
    -- CP-element group 1013: 	1020 
    -- CP-element group 1013:  members (1) 
      -- CP-element group 1013: 	 branch_block_stmt_714/ifx_xend1057_whilex_xbody898_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1013: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1013"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1006) & zeropad3D_CP_2152_elements(1009) & zeropad3D_CP_2152_elements(1012);
      gj_zeropad3D_cp_element_group_1013 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1013), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1014:  transition  output  delay-element  bypass 
    -- CP-element group 1014: predecessors 
    -- CP-element group 1014: 	446 
    -- CP-element group 1014: successors 
    -- CP-element group 1014: 	1019 
    -- CP-element group 1014:  members (4) 
      -- CP-element group 1014: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3154/$exit
      -- CP-element group 1014: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/$exit
      -- CP-element group 1014: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_sources/type_cast_3160_konst_delay_trans
      -- CP-element group 1014: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3154/phi_stmt_3154_req
      -- 
    phi_stmt_3154_req_13041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3154_req_13041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1014), ack => phi_stmt_3154_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1014) is a control-delay.
    cp_element_1014_delay: control_delay_element  generic map(name => " 1014_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(446), ack => zeropad3D_CP_2152_elements(1014), clk => clk, reset =>reset);
    -- CP-element group 1015:  transition  input  bypass 
    -- CP-element group 1015: predecessors 
    -- CP-element group 1015: 	446 
    -- CP-element group 1015: successors 
    -- CP-element group 1015: 	1017 
    -- CP-element group 1015:  members (2) 
      -- CP-element group 1015: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Sample/$exit
      -- CP-element group 1015: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Sample/ra
      -- 
    ra_13058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1015_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3151_inst_ack_0, ack => zeropad3D_CP_2152_elements(1015)); -- 
    -- CP-element group 1016:  transition  input  bypass 
    -- CP-element group 1016: predecessors 
    -- CP-element group 1016: 	446 
    -- CP-element group 1016: successors 
    -- CP-element group 1016: 	1017 
    -- CP-element group 1016:  members (2) 
      -- CP-element group 1016: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Update/$exit
      -- CP-element group 1016: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/Update/ca
      -- 
    ca_13063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1016_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3151_inst_ack_1, ack => zeropad3D_CP_2152_elements(1016)); -- 
    -- CP-element group 1017:  join  transition  output  bypass 
    -- CP-element group 1017: predecessors 
    -- CP-element group 1017: 	1015 
    -- CP-element group 1017: 	1016 
    -- CP-element group 1017: successors 
    -- CP-element group 1017: 	1019 
    -- CP-element group 1017:  members (5) 
      -- CP-element group 1017: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/$exit
      -- CP-element group 1017: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/$exit
      -- CP-element group 1017: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/$exit
      -- CP-element group 1017: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_sources/type_cast_3151/SplitProtocol/$exit
      -- CP-element group 1017: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3148/phi_stmt_3148_req
      -- 
    phi_stmt_3148_req_13064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3148_req_13064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1017), ack => phi_stmt_3148_req_0); -- 
    zeropad3D_cp_element_group_1017: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1017"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1015) & zeropad3D_CP_2152_elements(1016);
      gj_zeropad3D_cp_element_group_1017 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1017), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1018:  transition  output  delay-element  bypass 
    -- CP-element group 1018: predecessors 
    -- CP-element group 1018: 	446 
    -- CP-element group 1018: successors 
    -- CP-element group 1018: 	1019 
    -- CP-element group 1018:  members (4) 
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3141/$exit
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/$exit
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_sources/type_cast_3147_konst_delay_trans
      -- CP-element group 1018: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/phi_stmt_3141/phi_stmt_3141_req
      -- 
    phi_stmt_3141_req_13072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3141_req_13072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1018), ack => phi_stmt_3141_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1018) is a control-delay.
    cp_element_1018_delay: control_delay_element  generic map(name => " 1018_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(446), ack => zeropad3D_CP_2152_elements(1018), clk => clk, reset =>reset);
    -- CP-element group 1019:  join  transition  bypass 
    -- CP-element group 1019: predecessors 
    -- CP-element group 1019: 	1014 
    -- CP-element group 1019: 	1017 
    -- CP-element group 1019: 	1018 
    -- CP-element group 1019: successors 
    -- CP-element group 1019: 	1020 
    -- CP-element group 1019:  members (1) 
      -- CP-element group 1019: 	 branch_block_stmt_714/whilex_xend838_whilex_xbody898_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1019: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1019"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1014) & zeropad3D_CP_2152_elements(1017) & zeropad3D_CP_2152_elements(1018);
      gj_zeropad3D_cp_element_group_1019 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1019), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1020:  merge  fork  transition  place  bypass 
    -- CP-element group 1020: predecessors 
    -- CP-element group 1020: 	1013 
    -- CP-element group 1020: 	1019 
    -- CP-element group 1020: successors 
    -- CP-element group 1020: 	1021 
    -- CP-element group 1020: 	1022 
    -- CP-element group 1020: 	1023 
    -- CP-element group 1020:  members (2) 
      -- CP-element group 1020: 	 branch_block_stmt_714/merge_stmt_3140_PhiReqMerge
      -- CP-element group 1020: 	 branch_block_stmt_714/merge_stmt_3140_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1020) <= OrReduce(zeropad3D_CP_2152_elements(1013) & zeropad3D_CP_2152_elements(1019));
    -- CP-element group 1021:  transition  input  bypass 
    -- CP-element group 1021: predecessors 
    -- CP-element group 1021: 	1020 
    -- CP-element group 1021: successors 
    -- CP-element group 1021: 	1024 
    -- CP-element group 1021:  members (1) 
      -- CP-element group 1021: 	 branch_block_stmt_714/merge_stmt_3140_PhiAck/phi_stmt_3141_ack
      -- 
    phi_stmt_3141_ack_13077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1021_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3141_ack_0, ack => zeropad3D_CP_2152_elements(1021)); -- 
    -- CP-element group 1022:  transition  input  bypass 
    -- CP-element group 1022: predecessors 
    -- CP-element group 1022: 	1020 
    -- CP-element group 1022: successors 
    -- CP-element group 1022: 	1024 
    -- CP-element group 1022:  members (1) 
      -- CP-element group 1022: 	 branch_block_stmt_714/merge_stmt_3140_PhiAck/phi_stmt_3148_ack
      -- 
    phi_stmt_3148_ack_13078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1022_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3148_ack_0, ack => zeropad3D_CP_2152_elements(1022)); -- 
    -- CP-element group 1023:  transition  input  bypass 
    -- CP-element group 1023: predecessors 
    -- CP-element group 1023: 	1020 
    -- CP-element group 1023: successors 
    -- CP-element group 1023: 	1024 
    -- CP-element group 1023:  members (1) 
      -- CP-element group 1023: 	 branch_block_stmt_714/merge_stmt_3140_PhiAck/phi_stmt_3154_ack
      -- 
    phi_stmt_3154_ack_13079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1023_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3154_ack_0, ack => zeropad3D_CP_2152_elements(1023)); -- 
    -- CP-element group 1024:  join  fork  transition  place  output  bypass 
    -- CP-element group 1024: predecessors 
    -- CP-element group 1024: 	1021 
    -- CP-element group 1024: 	1022 
    -- CP-element group 1024: 	1023 
    -- CP-element group 1024: successors 
    -- CP-element group 1024: 	447 
    -- CP-element group 1024: 	448 
    -- CP-element group 1024:  members (10) 
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173__entry__
      -- CP-element group 1024: 	 branch_block_stmt_714/merge_stmt_3140__exit__
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/$entry
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_sample_start_
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_update_start_
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Sample/$entry
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Sample/rr
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Update/$entry
      -- CP-element group 1024: 	 branch_block_stmt_714/assign_stmt_3166_to_assign_stmt_3173/type_cast_3165_Update/cr
      -- CP-element group 1024: 	 branch_block_stmt_714/merge_stmt_3140_PhiAck/$exit
      -- 
    rr_7451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1024), ack => type_cast_3165_inst_req_0); -- 
    cr_7456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1024), ack => type_cast_3165_inst_req_1); -- 
    zeropad3D_cp_element_group_1024: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1024"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1021) & zeropad3D_CP_2152_elements(1022) & zeropad3D_CP_2152_elements(1023);
      gj_zeropad3D_cp_element_group_1024 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1024), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1025:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1025: predecessors 
    -- CP-element group 1025: 	449 
    -- CP-element group 1025: 	456 
    -- CP-element group 1025: 	459 
    -- CP-element group 1025: 	466 
    -- CP-element group 1025: successors 
    -- CP-element group 1025: 	467 
    -- CP-element group 1025: 	468 
    -- CP-element group 1025: 	469 
    -- CP-element group 1025: 	470 
    -- CP-element group 1025: 	473 
    -- CP-element group 1025: 	475 
    -- CP-element group 1025: 	477 
    -- CP-element group 1025: 	479 
    -- CP-element group 1025:  members (33) 
      -- CP-element group 1025: 	 branch_block_stmt_714/merge_stmt_3269__exit__
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325__entry__
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/word_access_complete/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/word_access_complete/word_0/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_Update/word_access_complete/word_0/cr
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_sample_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_update_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Sample/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Sample/rr
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Update/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3273_Update/cr
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_sample_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_update_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Sample/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Sample/rr
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Update/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3278_Update/cr
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_update_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Update/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/type_cast_3312_Update/cr
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_update_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_update_start
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Update/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/array_obj_ref_3318_final_index_sum_regn_Update/req
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_complete/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/addr_of_3319_complete/req
      -- CP-element group 1025: 	 branch_block_stmt_714/assign_stmt_3274_to_assign_stmt_3325/ptr_deref_3322_update_start_
      -- CP-element group 1025: 	 branch_block_stmt_714/merge_stmt_3269_PhiReqMerge
      -- CP-element group 1025: 	 branch_block_stmt_714/merge_stmt_3269_PhiAck/$entry
      -- CP-element group 1025: 	 branch_block_stmt_714/merge_stmt_3269_PhiAck/$exit
      -- CP-element group 1025: 	 branch_block_stmt_714/merge_stmt_3269_PhiAck/dummy
      -- 
    cr_7790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => ptr_deref_3322_store_0_req_1); -- 
    rr_7661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => type_cast_3273_inst_req_0); -- 
    cr_7666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => type_cast_3273_inst_req_1); -- 
    rr_7675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => type_cast_3278_inst_req_0); -- 
    cr_7680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => type_cast_3278_inst_req_1); -- 
    cr_7694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => type_cast_3312_inst_req_1); -- 
    req_7725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => array_obj_ref_3318_index_offset_req_1); -- 
    req_7740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1025), ack => addr_of_3319_final_reg_req_1); -- 
    zeropad3D_CP_2152_elements(1025) <= OrReduce(zeropad3D_CP_2152_elements(449) & zeropad3D_CP_2152_elements(456) & zeropad3D_CP_2152_elements(459) & zeropad3D_CP_2152_elements(466));
    -- CP-element group 1026:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1026: predecessors 
    -- CP-element group 1026: 	480 
    -- CP-element group 1026: 	500 
    -- CP-element group 1026: successors 
    -- CP-element group 1026: 	501 
    -- CP-element group 1026: 	502 
    -- CP-element group 1026:  members (13) 
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452__entry__
      -- CP-element group 1026: 	 branch_block_stmt_714/merge_stmt_3434__exit__
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/$entry
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_sample_start_
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_update_start_
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Sample/$entry
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Sample/rr
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Update/$entry
      -- CP-element group 1026: 	 branch_block_stmt_714/assign_stmt_3439_to_assign_stmt_3452/type_cast_3438_Update/cr
      -- CP-element group 1026: 	 branch_block_stmt_714/merge_stmt_3434_PhiReqMerge
      -- CP-element group 1026: 	 branch_block_stmt_714/merge_stmt_3434_PhiAck/$entry
      -- CP-element group 1026: 	 branch_block_stmt_714/merge_stmt_3434_PhiAck/$exit
      -- CP-element group 1026: 	 branch_block_stmt_714/merge_stmt_3434_PhiAck/dummy
      -- 
    rr_8039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1026), ack => type_cast_3438_inst_req_0); -- 
    cr_8044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1026), ack => type_cast_3438_inst_req_1); -- 
    zeropad3D_CP_2152_elements(1026) <= OrReduce(zeropad3D_CP_2152_elements(480) & zeropad3D_CP_2152_elements(500));
    -- CP-element group 1027:  transition  output  delay-element  bypass 
    -- CP-element group 1027: predecessors 
    -- CP-element group 1027: 	522 
    -- CP-element group 1027: successors 
    -- CP-element group 1027: 	1034 
    -- CP-element group 1027:  members (4) 
      -- CP-element group 1027: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3559/$exit
      -- CP-element group 1027: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/$exit
      -- CP-element group 1027: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3565_konst_delay_trans
      -- CP-element group 1027: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_req
      -- 
    phi_stmt_3559_req_13190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3559_req_13190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1027), ack => phi_stmt_3559_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1027) is a control-delay.
    cp_element_1027_delay: control_delay_element  generic map(name => " 1027_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(522), ack => zeropad3D_CP_2152_elements(1027), clk => clk, reset =>reset);
    -- CP-element group 1028:  transition  input  bypass 
    -- CP-element group 1028: predecessors 
    -- CP-element group 1028: 	522 
    -- CP-element group 1028: successors 
    -- CP-element group 1028: 	1030 
    -- CP-element group 1028:  members (2) 
      -- CP-element group 1028: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Sample/$exit
      -- CP-element group 1028: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Sample/ra
      -- 
    ra_13207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1028_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3571_inst_ack_0, ack => zeropad3D_CP_2152_elements(1028)); -- 
    -- CP-element group 1029:  transition  input  bypass 
    -- CP-element group 1029: predecessors 
    -- CP-element group 1029: 	522 
    -- CP-element group 1029: successors 
    -- CP-element group 1029: 	1030 
    -- CP-element group 1029:  members (2) 
      -- CP-element group 1029: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Update/$exit
      -- CP-element group 1029: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/Update/ca
      -- 
    ca_13212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1029_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3571_inst_ack_1, ack => zeropad3D_CP_2152_elements(1029)); -- 
    -- CP-element group 1030:  join  transition  output  bypass 
    -- CP-element group 1030: predecessors 
    -- CP-element group 1030: 	1028 
    -- CP-element group 1030: 	1029 
    -- CP-element group 1030: successors 
    -- CP-element group 1030: 	1034 
    -- CP-element group 1030:  members (5) 
      -- CP-element group 1030: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/$exit
      -- CP-element group 1030: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/$exit
      -- CP-element group 1030: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/$exit
      -- CP-element group 1030: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3571/SplitProtocol/$exit
      -- CP-element group 1030: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_req
      -- 
    phi_stmt_3566_req_13213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3566_req_13213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1030), ack => phi_stmt_3566_req_1); -- 
    zeropad3D_cp_element_group_1030: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1030"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1028) & zeropad3D_CP_2152_elements(1029);
      gj_zeropad3D_cp_element_group_1030 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1030), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1031:  transition  input  bypass 
    -- CP-element group 1031: predecessors 
    -- CP-element group 1031: 	522 
    -- CP-element group 1031: successors 
    -- CP-element group 1031: 	1033 
    -- CP-element group 1031:  members (2) 
      -- CP-element group 1031: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Sample/$exit
      -- CP-element group 1031: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Sample/ra
      -- 
    ra_13230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1031_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3575_inst_ack_0, ack => zeropad3D_CP_2152_elements(1031)); -- 
    -- CP-element group 1032:  transition  input  bypass 
    -- CP-element group 1032: predecessors 
    -- CP-element group 1032: 	522 
    -- CP-element group 1032: successors 
    -- CP-element group 1032: 	1033 
    -- CP-element group 1032:  members (2) 
      -- CP-element group 1032: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Update/$exit
      -- CP-element group 1032: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/Update/ca
      -- 
    ca_13235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1032_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3575_inst_ack_1, ack => zeropad3D_CP_2152_elements(1032)); -- 
    -- CP-element group 1033:  join  transition  output  bypass 
    -- CP-element group 1033: predecessors 
    -- CP-element group 1033: 	1031 
    -- CP-element group 1033: 	1032 
    -- CP-element group 1033: successors 
    -- CP-element group 1033: 	1034 
    -- CP-element group 1033:  members (5) 
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/$exit
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/$exit
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/$exit
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3575/SplitProtocol/$exit
      -- CP-element group 1033: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_req
      -- 
    phi_stmt_3572_req_13236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3572_req_13236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1033), ack => phi_stmt_3572_req_0); -- 
    zeropad3D_cp_element_group_1033: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1033"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1031) & zeropad3D_CP_2152_elements(1032);
      gj_zeropad3D_cp_element_group_1033 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1033), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1034:  join  transition  bypass 
    -- CP-element group 1034: predecessors 
    -- CP-element group 1034: 	1027 
    -- CP-element group 1034: 	1030 
    -- CP-element group 1034: 	1033 
    -- CP-element group 1034: successors 
    -- CP-element group 1034: 	1045 
    -- CP-element group 1034:  members (1) 
      -- CP-element group 1034: 	 branch_block_stmt_714/ifx_xelse1019_ifx_xend1057_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1034: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1034"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1027) & zeropad3D_CP_2152_elements(1030) & zeropad3D_CP_2152_elements(1033);
      gj_zeropad3D_cp_element_group_1034 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1034), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1035:  transition  input  bypass 
    -- CP-element group 1035: predecessors 
    -- CP-element group 1035: 	503 
    -- CP-element group 1035: successors 
    -- CP-element group 1035: 	1037 
    -- CP-element group 1035:  members (2) 
      -- CP-element group 1035: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Sample/$exit
      -- CP-element group 1035: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Sample/ra
      -- 
    ra_13256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1035_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3562_inst_ack_0, ack => zeropad3D_CP_2152_elements(1035)); -- 
    -- CP-element group 1036:  transition  input  bypass 
    -- CP-element group 1036: predecessors 
    -- CP-element group 1036: 	503 
    -- CP-element group 1036: successors 
    -- CP-element group 1036: 	1037 
    -- CP-element group 1036:  members (2) 
      -- CP-element group 1036: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Update/$exit
      -- CP-element group 1036: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/Update/ca
      -- 
    ca_13261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1036_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3562_inst_ack_1, ack => zeropad3D_CP_2152_elements(1036)); -- 
    -- CP-element group 1037:  join  transition  output  bypass 
    -- CP-element group 1037: predecessors 
    -- CP-element group 1037: 	1035 
    -- CP-element group 1037: 	1036 
    -- CP-element group 1037: successors 
    -- CP-element group 1037: 	1044 
    -- CP-element group 1037:  members (5) 
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_sources/type_cast_3562/SplitProtocol/$exit
      -- CP-element group 1037: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3559/phi_stmt_3559_req
      -- 
    phi_stmt_3559_req_13262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3559_req_13262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1037), ack => phi_stmt_3559_req_0); -- 
    zeropad3D_cp_element_group_1037: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1037"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1035) & zeropad3D_CP_2152_elements(1036);
      gj_zeropad3D_cp_element_group_1037 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1037), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1038:  transition  input  bypass 
    -- CP-element group 1038: predecessors 
    -- CP-element group 1038: 	503 
    -- CP-element group 1038: successors 
    -- CP-element group 1038: 	1040 
    -- CP-element group 1038:  members (2) 
      -- CP-element group 1038: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Sample/$exit
      -- CP-element group 1038: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Sample/ra
      -- 
    ra_13279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1038_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3569_inst_ack_0, ack => zeropad3D_CP_2152_elements(1038)); -- 
    -- CP-element group 1039:  transition  input  bypass 
    -- CP-element group 1039: predecessors 
    -- CP-element group 1039: 	503 
    -- CP-element group 1039: successors 
    -- CP-element group 1039: 	1040 
    -- CP-element group 1039:  members (2) 
      -- CP-element group 1039: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Update/$exit
      -- CP-element group 1039: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/Update/ca
      -- 
    ca_13284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1039_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3569_inst_ack_1, ack => zeropad3D_CP_2152_elements(1039)); -- 
    -- CP-element group 1040:  join  transition  output  bypass 
    -- CP-element group 1040: predecessors 
    -- CP-element group 1040: 	1038 
    -- CP-element group 1040: 	1039 
    -- CP-element group 1040: successors 
    -- CP-element group 1040: 	1044 
    -- CP-element group 1040:  members (5) 
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/$exit
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/$exit
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/$exit
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_sources/type_cast_3569/SplitProtocol/$exit
      -- CP-element group 1040: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3566/phi_stmt_3566_req
      -- 
    phi_stmt_3566_req_13285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3566_req_13285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1040), ack => phi_stmt_3566_req_0); -- 
    zeropad3D_cp_element_group_1040: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1040"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1038) & zeropad3D_CP_2152_elements(1039);
      gj_zeropad3D_cp_element_group_1040 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1040), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1041:  transition  input  bypass 
    -- CP-element group 1041: predecessors 
    -- CP-element group 1041: 	503 
    -- CP-element group 1041: successors 
    -- CP-element group 1041: 	1043 
    -- CP-element group 1041:  members (2) 
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Sample/$exit
      -- CP-element group 1041: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Sample/ra
      -- 
    ra_13302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1041_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3577_inst_ack_0, ack => zeropad3D_CP_2152_elements(1041)); -- 
    -- CP-element group 1042:  transition  input  bypass 
    -- CP-element group 1042: predecessors 
    -- CP-element group 1042: 	503 
    -- CP-element group 1042: successors 
    -- CP-element group 1042: 	1043 
    -- CP-element group 1042:  members (2) 
      -- CP-element group 1042: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Update/$exit
      -- CP-element group 1042: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/Update/ca
      -- 
    ca_13307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1042_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3577_inst_ack_1, ack => zeropad3D_CP_2152_elements(1042)); -- 
    -- CP-element group 1043:  join  transition  output  bypass 
    -- CP-element group 1043: predecessors 
    -- CP-element group 1043: 	1041 
    -- CP-element group 1043: 	1042 
    -- CP-element group 1043: successors 
    -- CP-element group 1043: 	1044 
    -- CP-element group 1043:  members (5) 
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/$exit
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/$exit
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/$exit
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_sources/type_cast_3577/SplitProtocol/$exit
      -- CP-element group 1043: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/phi_stmt_3572/phi_stmt_3572_req
      -- 
    phi_stmt_3572_req_13308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3572_req_13308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1043), ack => phi_stmt_3572_req_1); -- 
    zeropad3D_cp_element_group_1043: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1043"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1041) & zeropad3D_CP_2152_elements(1042);
      gj_zeropad3D_cp_element_group_1043 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1043), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1044:  join  transition  bypass 
    -- CP-element group 1044: predecessors 
    -- CP-element group 1044: 	1037 
    -- CP-element group 1044: 	1040 
    -- CP-element group 1044: 	1043 
    -- CP-element group 1044: successors 
    -- CP-element group 1044: 	1045 
    -- CP-element group 1044:  members (1) 
      -- CP-element group 1044: 	 branch_block_stmt_714/ifx_xthen1014_ifx_xend1057_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1044: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1044"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1037) & zeropad3D_CP_2152_elements(1040) & zeropad3D_CP_2152_elements(1043);
      gj_zeropad3D_cp_element_group_1044 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1044), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1045:  merge  fork  transition  place  bypass 
    -- CP-element group 1045: predecessors 
    -- CP-element group 1045: 	1034 
    -- CP-element group 1045: 	1044 
    -- CP-element group 1045: successors 
    -- CP-element group 1045: 	1046 
    -- CP-element group 1045: 	1047 
    -- CP-element group 1045: 	1048 
    -- CP-element group 1045:  members (2) 
      -- CP-element group 1045: 	 branch_block_stmt_714/merge_stmt_3558_PhiReqMerge
      -- CP-element group 1045: 	 branch_block_stmt_714/merge_stmt_3558_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1045) <= OrReduce(zeropad3D_CP_2152_elements(1034) & zeropad3D_CP_2152_elements(1044));
    -- CP-element group 1046:  transition  input  bypass 
    -- CP-element group 1046: predecessors 
    -- CP-element group 1046: 	1045 
    -- CP-element group 1046: successors 
    -- CP-element group 1046: 	1049 
    -- CP-element group 1046:  members (1) 
      -- CP-element group 1046: 	 branch_block_stmt_714/merge_stmt_3558_PhiAck/phi_stmt_3559_ack
      -- 
    phi_stmt_3559_ack_13313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1046_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3559_ack_0, ack => zeropad3D_CP_2152_elements(1046)); -- 
    -- CP-element group 1047:  transition  input  bypass 
    -- CP-element group 1047: predecessors 
    -- CP-element group 1047: 	1045 
    -- CP-element group 1047: successors 
    -- CP-element group 1047: 	1049 
    -- CP-element group 1047:  members (1) 
      -- CP-element group 1047: 	 branch_block_stmt_714/merge_stmt_3558_PhiAck/phi_stmt_3566_ack
      -- 
    phi_stmt_3566_ack_13314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1047_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3566_ack_0, ack => zeropad3D_CP_2152_elements(1047)); -- 
    -- CP-element group 1048:  transition  input  bypass 
    -- CP-element group 1048: predecessors 
    -- CP-element group 1048: 	1045 
    -- CP-element group 1048: successors 
    -- CP-element group 1048: 	1049 
    -- CP-element group 1048:  members (1) 
      -- CP-element group 1048: 	 branch_block_stmt_714/merge_stmt_3558_PhiAck/phi_stmt_3572_ack
      -- 
    phi_stmt_3572_ack_13315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1048_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3572_ack_0, ack => zeropad3D_CP_2152_elements(1048)); -- 
    -- CP-element group 1049:  join  transition  bypass 
    -- CP-element group 1049: predecessors 
    -- CP-element group 1049: 	1046 
    -- CP-element group 1049: 	1047 
    -- CP-element group 1049: 	1048 
    -- CP-element group 1049: successors 
    -- CP-element group 1049: 	5 
    -- CP-element group 1049:  members (1) 
      -- CP-element group 1049: 	 branch_block_stmt_714/merge_stmt_3558_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1049: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1049"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1046) & zeropad3D_CP_2152_elements(1047) & zeropad3D_CP_2152_elements(1048);
      gj_zeropad3D_cp_element_group_1049 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1049), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1050:  transition  input  bypass 
    -- CP-element group 1050: predecessors 
    -- CP-element group 1050: 	6 
    -- CP-element group 1050: successors 
    -- CP-element group 1050: 	1052 
    -- CP-element group 1050:  members (2) 
      -- CP-element group 1050: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/$exit
      -- CP-element group 1050: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Sample/ra
      -- 
    ra_13343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1050_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3731_inst_ack_0, ack => zeropad3D_CP_2152_elements(1050)); -- 
    -- CP-element group 1051:  transition  input  bypass 
    -- CP-element group 1051: predecessors 
    -- CP-element group 1051: 	6 
    -- CP-element group 1051: successors 
    -- CP-element group 1051: 	1052 
    -- CP-element group 1051:  members (2) 
      -- CP-element group 1051: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/$exit
      -- CP-element group 1051: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/Update/ca
      -- 
    ca_13348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1051_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3731_inst_ack_1, ack => zeropad3D_CP_2152_elements(1051)); -- 
    -- CP-element group 1052:  join  transition  output  bypass 
    -- CP-element group 1052: predecessors 
    -- CP-element group 1052: 	1050 
    -- CP-element group 1052: 	1051 
    -- CP-element group 1052: successors 
    -- CP-element group 1052: 	1059 
    -- CP-element group 1052:  members (5) 
      -- CP-element group 1052: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/$exit
      -- CP-element group 1052: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$exit
      -- CP-element group 1052: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/$exit
      -- CP-element group 1052: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3731/SplitProtocol/$exit
      -- CP-element group 1052: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_req
      -- 
    phi_stmt_3728_req_13349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3728_req_13349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1052), ack => phi_stmt_3728_req_0); -- 
    zeropad3D_cp_element_group_1052: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1052"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1050) & zeropad3D_CP_2152_elements(1051);
      gj_zeropad3D_cp_element_group_1052 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1052), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1053:  transition  input  bypass 
    -- CP-element group 1053: predecessors 
    -- CP-element group 1053: 	6 
    -- CP-element group 1053: successors 
    -- CP-element group 1053: 	1055 
    -- CP-element group 1053:  members (2) 
      -- CP-element group 1053: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Sample/$exit
      -- CP-element group 1053: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Sample/ra
      -- 
    ra_13366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1053_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3740_inst_ack_0, ack => zeropad3D_CP_2152_elements(1053)); -- 
    -- CP-element group 1054:  transition  input  bypass 
    -- CP-element group 1054: predecessors 
    -- CP-element group 1054: 	6 
    -- CP-element group 1054: successors 
    -- CP-element group 1054: 	1055 
    -- CP-element group 1054:  members (2) 
      -- CP-element group 1054: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Update/$exit
      -- CP-element group 1054: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/Update/ca
      -- 
    ca_13371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1054_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3740_inst_ack_1, ack => zeropad3D_CP_2152_elements(1054)); -- 
    -- CP-element group 1055:  join  transition  output  bypass 
    -- CP-element group 1055: predecessors 
    -- CP-element group 1055: 	1053 
    -- CP-element group 1055: 	1054 
    -- CP-element group 1055: successors 
    -- CP-element group 1055: 	1059 
    -- CP-element group 1055:  members (5) 
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/$exit
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/$exit
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/$exit
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3740/SplitProtocol/$exit
      -- CP-element group 1055: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_req
      -- 
    phi_stmt_3735_req_13372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3735_req_13372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1055), ack => phi_stmt_3735_req_1); -- 
    zeropad3D_cp_element_group_1055: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1055"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1053) & zeropad3D_CP_2152_elements(1054);
      gj_zeropad3D_cp_element_group_1055 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1055), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1056:  transition  input  bypass 
    -- CP-element group 1056: predecessors 
    -- CP-element group 1056: 	6 
    -- CP-element group 1056: successors 
    -- CP-element group 1056: 	1058 
    -- CP-element group 1056:  members (2) 
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Sample/$exit
      -- CP-element group 1056: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Sample/ra
      -- 
    ra_13389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1056_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3744_inst_ack_0, ack => zeropad3D_CP_2152_elements(1056)); -- 
    -- CP-element group 1057:  transition  input  bypass 
    -- CP-element group 1057: predecessors 
    -- CP-element group 1057: 	6 
    -- CP-element group 1057: successors 
    -- CP-element group 1057: 	1058 
    -- CP-element group 1057:  members (2) 
      -- CP-element group 1057: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Update/$exit
      -- CP-element group 1057: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/Update/ca
      -- 
    ca_13394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1057_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3744_inst_ack_1, ack => zeropad3D_CP_2152_elements(1057)); -- 
    -- CP-element group 1058:  join  transition  output  bypass 
    -- CP-element group 1058: predecessors 
    -- CP-element group 1058: 	1056 
    -- CP-element group 1058: 	1057 
    -- CP-element group 1058: successors 
    -- CP-element group 1058: 	1059 
    -- CP-element group 1058:  members (5) 
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/$exit
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/$exit
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/$exit
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3744/SplitProtocol/$exit
      -- CP-element group 1058: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_req
      -- 
    phi_stmt_3741_req_13395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3741_req_13395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1058), ack => phi_stmt_3741_req_0); -- 
    zeropad3D_cp_element_group_1058: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1058"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1056) & zeropad3D_CP_2152_elements(1057);
      gj_zeropad3D_cp_element_group_1058 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1058), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1059:  join  transition  bypass 
    -- CP-element group 1059: predecessors 
    -- CP-element group 1059: 	1052 
    -- CP-element group 1059: 	1055 
    -- CP-element group 1059: 	1058 
    -- CP-element group 1059: successors 
    -- CP-element group 1059: 	1068 
    -- CP-element group 1059:  members (1) 
      -- CP-element group 1059: 	 branch_block_stmt_714/ifx_xend1279_whilex_xbody1122_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1059: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1059"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1052) & zeropad3D_CP_2152_elements(1055) & zeropad3D_CP_2152_elements(1058);
      gj_zeropad3D_cp_element_group_1059 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1059), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1060:  transition  output  delay-element  bypass 
    -- CP-element group 1060: predecessors 
    -- CP-element group 1060: 	545 
    -- CP-element group 1060: successors 
    -- CP-element group 1060: 	1067 
    -- CP-element group 1060:  members (4) 
      -- CP-element group 1060: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3728/$exit
      -- CP-element group 1060: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/$exit
      -- CP-element group 1060: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_sources/type_cast_3734_konst_delay_trans
      -- CP-element group 1060: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3728/phi_stmt_3728_req
      -- 
    phi_stmt_3728_req_13406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3728_req_13406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1060), ack => phi_stmt_3728_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1060) is a control-delay.
    cp_element_1060_delay: control_delay_element  generic map(name => " 1060_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(545), ack => zeropad3D_CP_2152_elements(1060), clk => clk, reset =>reset);
    -- CP-element group 1061:  transition  input  bypass 
    -- CP-element group 1061: predecessors 
    -- CP-element group 1061: 	545 
    -- CP-element group 1061: successors 
    -- CP-element group 1061: 	1063 
    -- CP-element group 1061:  members (2) 
      -- CP-element group 1061: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Sample/$exit
      -- CP-element group 1061: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Sample/ra
      -- 
    ra_13423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1061_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3738_inst_ack_0, ack => zeropad3D_CP_2152_elements(1061)); -- 
    -- CP-element group 1062:  transition  input  bypass 
    -- CP-element group 1062: predecessors 
    -- CP-element group 1062: 	545 
    -- CP-element group 1062: successors 
    -- CP-element group 1062: 	1063 
    -- CP-element group 1062:  members (2) 
      -- CP-element group 1062: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Update/$exit
      -- CP-element group 1062: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/Update/ca
      -- 
    ca_13428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1062_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3738_inst_ack_1, ack => zeropad3D_CP_2152_elements(1062)); -- 
    -- CP-element group 1063:  join  transition  output  bypass 
    -- CP-element group 1063: predecessors 
    -- CP-element group 1063: 	1061 
    -- CP-element group 1063: 	1062 
    -- CP-element group 1063: successors 
    -- CP-element group 1063: 	1067 
    -- CP-element group 1063:  members (5) 
      -- CP-element group 1063: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/$exit
      -- CP-element group 1063: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/$exit
      -- CP-element group 1063: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/$exit
      -- CP-element group 1063: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_sources/type_cast_3738/SplitProtocol/$exit
      -- CP-element group 1063: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3735/phi_stmt_3735_req
      -- 
    phi_stmt_3735_req_13429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3735_req_13429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1063), ack => phi_stmt_3735_req_0); -- 
    zeropad3D_cp_element_group_1063: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1063"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1061) & zeropad3D_CP_2152_elements(1062);
      gj_zeropad3D_cp_element_group_1063 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1063), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1064:  transition  input  bypass 
    -- CP-element group 1064: predecessors 
    -- CP-element group 1064: 	545 
    -- CP-element group 1064: successors 
    -- CP-element group 1064: 	1066 
    -- CP-element group 1064:  members (2) 
      -- CP-element group 1064: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Sample/$exit
      -- CP-element group 1064: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Sample/ra
      -- 
    ra_13446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1064_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3746_inst_ack_0, ack => zeropad3D_CP_2152_elements(1064)); -- 
    -- CP-element group 1065:  transition  input  bypass 
    -- CP-element group 1065: predecessors 
    -- CP-element group 1065: 	545 
    -- CP-element group 1065: successors 
    -- CP-element group 1065: 	1066 
    -- CP-element group 1065:  members (2) 
      -- CP-element group 1065: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Update/$exit
      -- CP-element group 1065: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/Update/ca
      -- 
    ca_13451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1065_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3746_inst_ack_1, ack => zeropad3D_CP_2152_elements(1065)); -- 
    -- CP-element group 1066:  join  transition  output  bypass 
    -- CP-element group 1066: predecessors 
    -- CP-element group 1066: 	1064 
    -- CP-element group 1066: 	1065 
    -- CP-element group 1066: successors 
    -- CP-element group 1066: 	1067 
    -- CP-element group 1066:  members (5) 
      -- CP-element group 1066: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/$exit
      -- CP-element group 1066: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/$exit
      -- CP-element group 1066: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/$exit
      -- CP-element group 1066: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_sources/type_cast_3746/SplitProtocol/$exit
      -- CP-element group 1066: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/phi_stmt_3741/phi_stmt_3741_req
      -- 
    phi_stmt_3741_req_13452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3741_req_13452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1066), ack => phi_stmt_3741_req_1); -- 
    zeropad3D_cp_element_group_1066: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1066"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1064) & zeropad3D_CP_2152_elements(1065);
      gj_zeropad3D_cp_element_group_1066 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1066), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1067:  join  transition  bypass 
    -- CP-element group 1067: predecessors 
    -- CP-element group 1067: 	1060 
    -- CP-element group 1067: 	1063 
    -- CP-element group 1067: 	1066 
    -- CP-element group 1067: successors 
    -- CP-element group 1067: 	1068 
    -- CP-element group 1067:  members (1) 
      -- CP-element group 1067: 	 branch_block_stmt_714/whilex_xend1058_whilex_xbody1122_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1067: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1067"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1060) & zeropad3D_CP_2152_elements(1063) & zeropad3D_CP_2152_elements(1066);
      gj_zeropad3D_cp_element_group_1067 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1067), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1068:  merge  fork  transition  place  bypass 
    -- CP-element group 1068: predecessors 
    -- CP-element group 1068: 	1059 
    -- CP-element group 1068: 	1067 
    -- CP-element group 1068: successors 
    -- CP-element group 1068: 	1069 
    -- CP-element group 1068: 	1070 
    -- CP-element group 1068: 	1071 
    -- CP-element group 1068:  members (2) 
      -- CP-element group 1068: 	 branch_block_stmt_714/merge_stmt_3727_PhiReqMerge
      -- CP-element group 1068: 	 branch_block_stmt_714/merge_stmt_3727_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1068) <= OrReduce(zeropad3D_CP_2152_elements(1059) & zeropad3D_CP_2152_elements(1067));
    -- CP-element group 1069:  transition  input  bypass 
    -- CP-element group 1069: predecessors 
    -- CP-element group 1069: 	1068 
    -- CP-element group 1069: successors 
    -- CP-element group 1069: 	1072 
    -- CP-element group 1069:  members (1) 
      -- CP-element group 1069: 	 branch_block_stmt_714/merge_stmt_3727_PhiAck/phi_stmt_3728_ack
      -- 
    phi_stmt_3728_ack_13457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1069_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3728_ack_0, ack => zeropad3D_CP_2152_elements(1069)); -- 
    -- CP-element group 1070:  transition  input  bypass 
    -- CP-element group 1070: predecessors 
    -- CP-element group 1070: 	1068 
    -- CP-element group 1070: successors 
    -- CP-element group 1070: 	1072 
    -- CP-element group 1070:  members (1) 
      -- CP-element group 1070: 	 branch_block_stmt_714/merge_stmt_3727_PhiAck/phi_stmt_3735_ack
      -- 
    phi_stmt_3735_ack_13458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1070_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3735_ack_0, ack => zeropad3D_CP_2152_elements(1070)); -- 
    -- CP-element group 1071:  transition  input  bypass 
    -- CP-element group 1071: predecessors 
    -- CP-element group 1071: 	1068 
    -- CP-element group 1071: successors 
    -- CP-element group 1071: 	1072 
    -- CP-element group 1071:  members (1) 
      -- CP-element group 1071: 	 branch_block_stmt_714/merge_stmt_3727_PhiAck/phi_stmt_3741_ack
      -- 
    phi_stmt_3741_ack_13459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1071_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3741_ack_0, ack => zeropad3D_CP_2152_elements(1071)); -- 
    -- CP-element group 1072:  join  fork  transition  place  output  bypass 
    -- CP-element group 1072: predecessors 
    -- CP-element group 1072: 	1069 
    -- CP-element group 1072: 	1070 
    -- CP-element group 1072: 	1071 
    -- CP-element group 1072: successors 
    -- CP-element group 1072: 	546 
    -- CP-element group 1072: 	547 
    -- CP-element group 1072:  members (10) 
      -- CP-element group 1072: 	 branch_block_stmt_714/merge_stmt_3727__exit__
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759__entry__
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/$entry
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_sample_start_
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_update_start_
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Sample/$entry
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Sample/rr
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Update/$entry
      -- CP-element group 1072: 	 branch_block_stmt_714/assign_stmt_3752_to_assign_stmt_3759/type_cast_3751_Update/cr
      -- CP-element group 1072: 	 branch_block_stmt_714/merge_stmt_3727_PhiAck/$exit
      -- 
    rr_8541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1072), ack => type_cast_3751_inst_req_0); -- 
    cr_8546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1072), ack => type_cast_3751_inst_req_1); -- 
    zeropad3D_cp_element_group_1072: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1072"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1069) & zeropad3D_CP_2152_elements(1070) & zeropad3D_CP_2152_elements(1071);
      gj_zeropad3D_cp_element_group_1072 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1072), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1073:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1073: predecessors 
    -- CP-element group 1073: 	548 
    -- CP-element group 1073: 	555 
    -- CP-element group 1073: 	558 
    -- CP-element group 1073: 	565 
    -- CP-element group 1073: successors 
    -- CP-element group 1073: 	566 
    -- CP-element group 1073: 	567 
    -- CP-element group 1073: 	568 
    -- CP-element group 1073: 	569 
    -- CP-element group 1073: 	572 
    -- CP-element group 1073: 	574 
    -- CP-element group 1073: 	576 
    -- CP-element group 1073: 	578 
    -- CP-element group 1073:  members (33) 
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905__entry__
      -- CP-element group 1073: 	 branch_block_stmt_714/merge_stmt_3849__exit__
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_sample_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_update_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Sample/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Sample/rr
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Update/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3853_Update/cr
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_sample_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_update_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Sample/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Sample/rr
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Update/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3858_Update/cr
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_update_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Update/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/type_cast_3892_Update/cr
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_update_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_update_start
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Update/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/array_obj_ref_3898_final_index_sum_regn_Update/req
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_complete/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/addr_of_3899_complete/req
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_update_start_
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/word_access_complete/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/word_access_complete/word_0/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/assign_stmt_3854_to_assign_stmt_3905/ptr_deref_3902_Update/word_access_complete/word_0/cr
      -- CP-element group 1073: 	 branch_block_stmt_714/merge_stmt_3849_PhiReqMerge
      -- CP-element group 1073: 	 branch_block_stmt_714/merge_stmt_3849_PhiAck/$entry
      -- CP-element group 1073: 	 branch_block_stmt_714/merge_stmt_3849_PhiAck/$exit
      -- CP-element group 1073: 	 branch_block_stmt_714/merge_stmt_3849_PhiAck/dummy
      -- 
    rr_8751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => type_cast_3853_inst_req_0); -- 
    cr_8756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => type_cast_3853_inst_req_1); -- 
    rr_8765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => type_cast_3858_inst_req_0); -- 
    cr_8770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => type_cast_3858_inst_req_1); -- 
    cr_8784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => type_cast_3892_inst_req_1); -- 
    req_8815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => array_obj_ref_3898_index_offset_req_1); -- 
    req_8830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => addr_of_3899_final_reg_req_1); -- 
    cr_8880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1073), ack => ptr_deref_3902_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(1073) <= OrReduce(zeropad3D_CP_2152_elements(548) & zeropad3D_CP_2152_elements(555) & zeropad3D_CP_2152_elements(558) & zeropad3D_CP_2152_elements(565));
    -- CP-element group 1074:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1074: predecessors 
    -- CP-element group 1074: 	579 
    -- CP-element group 1074: 	599 
    -- CP-element group 1074: successors 
    -- CP-element group 1074: 	600 
    -- CP-element group 1074: 	601 
    -- CP-element group 1074:  members (13) 
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032__entry__
      -- CP-element group 1074: 	 branch_block_stmt_714/merge_stmt_4014__exit__
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/$entry
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_sample_start_
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_update_start_
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Sample/$entry
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Sample/rr
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Update/$entry
      -- CP-element group 1074: 	 branch_block_stmt_714/assign_stmt_4019_to_assign_stmt_4032/type_cast_4018_Update/cr
      -- CP-element group 1074: 	 branch_block_stmt_714/merge_stmt_4014_PhiReqMerge
      -- CP-element group 1074: 	 branch_block_stmt_714/merge_stmt_4014_PhiAck/$entry
      -- CP-element group 1074: 	 branch_block_stmt_714/merge_stmt_4014_PhiAck/$exit
      -- CP-element group 1074: 	 branch_block_stmt_714/merge_stmt_4014_PhiAck/dummy
      -- 
    rr_9129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1074), ack => type_cast_4018_inst_req_0); -- 
    cr_9134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1074), ack => type_cast_4018_inst_req_1); -- 
    zeropad3D_CP_2152_elements(1074) <= OrReduce(zeropad3D_CP_2152_elements(579) & zeropad3D_CP_2152_elements(599));
    -- CP-element group 1075:  transition  output  delay-element  bypass 
    -- CP-element group 1075: predecessors 
    -- CP-element group 1075: 	621 
    -- CP-element group 1075: successors 
    -- CP-element group 1075: 	1082 
    -- CP-element group 1075:  members (4) 
      -- CP-element group 1075: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4132/$exit
      -- CP-element group 1075: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/$exit
      -- CP-element group 1075: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4138_konst_delay_trans
      -- CP-element group 1075: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_req
      -- 
    phi_stmt_4132_req_13570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4132_req_13570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1075), ack => phi_stmt_4132_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1075) is a control-delay.
    cp_element_1075_delay: control_delay_element  generic map(name => " 1075_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(621), ack => zeropad3D_CP_2152_elements(1075), clk => clk, reset =>reset);
    -- CP-element group 1076:  transition  input  bypass 
    -- CP-element group 1076: predecessors 
    -- CP-element group 1076: 	621 
    -- CP-element group 1076: successors 
    -- CP-element group 1076: 	1078 
    -- CP-element group 1076:  members (2) 
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Sample/$exit
      -- CP-element group 1076: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Sample/ra
      -- 
    ra_13587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1076_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4144_inst_ack_0, ack => zeropad3D_CP_2152_elements(1076)); -- 
    -- CP-element group 1077:  transition  input  bypass 
    -- CP-element group 1077: predecessors 
    -- CP-element group 1077: 	621 
    -- CP-element group 1077: successors 
    -- CP-element group 1077: 	1078 
    -- CP-element group 1077:  members (2) 
      -- CP-element group 1077: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Update/$exit
      -- CP-element group 1077: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/Update/ca
      -- 
    ca_13592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1077_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4144_inst_ack_1, ack => zeropad3D_CP_2152_elements(1077)); -- 
    -- CP-element group 1078:  join  transition  output  bypass 
    -- CP-element group 1078: predecessors 
    -- CP-element group 1078: 	1076 
    -- CP-element group 1078: 	1077 
    -- CP-element group 1078: successors 
    -- CP-element group 1078: 	1082 
    -- CP-element group 1078:  members (5) 
      -- CP-element group 1078: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/$exit
      -- CP-element group 1078: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/$exit
      -- CP-element group 1078: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/$exit
      -- CP-element group 1078: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4144/SplitProtocol/$exit
      -- CP-element group 1078: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_req
      -- 
    phi_stmt_4139_req_13593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4139_req_13593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1078), ack => phi_stmt_4139_req_1); -- 
    zeropad3D_cp_element_group_1078: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1078"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1076) & zeropad3D_CP_2152_elements(1077);
      gj_zeropad3D_cp_element_group_1078 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1078), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1079:  transition  input  bypass 
    -- CP-element group 1079: predecessors 
    -- CP-element group 1079: 	621 
    -- CP-element group 1079: successors 
    -- CP-element group 1079: 	1081 
    -- CP-element group 1079:  members (2) 
      -- CP-element group 1079: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Sample/$exit
      -- CP-element group 1079: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Sample/ra
      -- 
    ra_13610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1079_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4150_inst_ack_0, ack => zeropad3D_CP_2152_elements(1079)); -- 
    -- CP-element group 1080:  transition  input  bypass 
    -- CP-element group 1080: predecessors 
    -- CP-element group 1080: 	621 
    -- CP-element group 1080: successors 
    -- CP-element group 1080: 	1081 
    -- CP-element group 1080:  members (2) 
      -- CP-element group 1080: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Update/$exit
      -- CP-element group 1080: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/Update/ca
      -- 
    ca_13615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1080_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4150_inst_ack_1, ack => zeropad3D_CP_2152_elements(1080)); -- 
    -- CP-element group 1081:  join  transition  output  bypass 
    -- CP-element group 1081: predecessors 
    -- CP-element group 1081: 	1079 
    -- CP-element group 1081: 	1080 
    -- CP-element group 1081: successors 
    -- CP-element group 1081: 	1082 
    -- CP-element group 1081:  members (5) 
      -- CP-element group 1081: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4150/SplitProtocol/$exit
      -- CP-element group 1081: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_req
      -- 
    phi_stmt_4145_req_13616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4145_req_13616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1081), ack => phi_stmt_4145_req_1); -- 
    zeropad3D_cp_element_group_1081: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1081"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1079) & zeropad3D_CP_2152_elements(1080);
      gj_zeropad3D_cp_element_group_1081 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1081), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1082:  join  transition  bypass 
    -- CP-element group 1082: predecessors 
    -- CP-element group 1082: 	1075 
    -- CP-element group 1082: 	1078 
    -- CP-element group 1082: 	1081 
    -- CP-element group 1082: successors 
    -- CP-element group 1082: 	1093 
    -- CP-element group 1082:  members (1) 
      -- CP-element group 1082: 	 branch_block_stmt_714/ifx_xelse1242_ifx_xend1279_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1082: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1082"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1075) & zeropad3D_CP_2152_elements(1078) & zeropad3D_CP_2152_elements(1081);
      gj_zeropad3D_cp_element_group_1082 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1082), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1083:  transition  input  bypass 
    -- CP-element group 1083: predecessors 
    -- CP-element group 1083: 	602 
    -- CP-element group 1083: successors 
    -- CP-element group 1083: 	1085 
    -- CP-element group 1083:  members (2) 
      -- CP-element group 1083: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Sample/$exit
      -- CP-element group 1083: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Sample/ra
      -- 
    ra_13636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1083_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4135_inst_ack_0, ack => zeropad3D_CP_2152_elements(1083)); -- 
    -- CP-element group 1084:  transition  input  bypass 
    -- CP-element group 1084: predecessors 
    -- CP-element group 1084: 	602 
    -- CP-element group 1084: successors 
    -- CP-element group 1084: 	1085 
    -- CP-element group 1084:  members (2) 
      -- CP-element group 1084: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Update/$exit
      -- CP-element group 1084: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/Update/ca
      -- 
    ca_13641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1084_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4135_inst_ack_1, ack => zeropad3D_CP_2152_elements(1084)); -- 
    -- CP-element group 1085:  join  transition  output  bypass 
    -- CP-element group 1085: predecessors 
    -- CP-element group 1085: 	1083 
    -- CP-element group 1085: 	1084 
    -- CP-element group 1085: successors 
    -- CP-element group 1085: 	1092 
    -- CP-element group 1085:  members (5) 
      -- CP-element group 1085: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/$exit
      -- CP-element group 1085: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/$exit
      -- CP-element group 1085: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/$exit
      -- CP-element group 1085: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_sources/type_cast_4135/SplitProtocol/$exit
      -- CP-element group 1085: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4132/phi_stmt_4132_req
      -- 
    phi_stmt_4132_req_13642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4132_req_13642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1085), ack => phi_stmt_4132_req_0); -- 
    zeropad3D_cp_element_group_1085: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1085"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1083) & zeropad3D_CP_2152_elements(1084);
      gj_zeropad3D_cp_element_group_1085 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1085), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1086:  transition  input  bypass 
    -- CP-element group 1086: predecessors 
    -- CP-element group 1086: 	602 
    -- CP-element group 1086: successors 
    -- CP-element group 1086: 	1088 
    -- CP-element group 1086:  members (2) 
      -- CP-element group 1086: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Sample/ra
      -- CP-element group 1086: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Sample/$exit
      -- 
    ra_13659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1086_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4142_inst_ack_0, ack => zeropad3D_CP_2152_elements(1086)); -- 
    -- CP-element group 1087:  transition  input  bypass 
    -- CP-element group 1087: predecessors 
    -- CP-element group 1087: 	602 
    -- CP-element group 1087: successors 
    -- CP-element group 1087: 	1088 
    -- CP-element group 1087:  members (2) 
      -- CP-element group 1087: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Update/ca
      -- CP-element group 1087: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/Update/$exit
      -- 
    ca_13664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1087_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4142_inst_ack_1, ack => zeropad3D_CP_2152_elements(1087)); -- 
    -- CP-element group 1088:  join  transition  output  bypass 
    -- CP-element group 1088: predecessors 
    -- CP-element group 1088: 	1086 
    -- CP-element group 1088: 	1087 
    -- CP-element group 1088: successors 
    -- CP-element group 1088: 	1092 
    -- CP-element group 1088:  members (5) 
      -- CP-element group 1088: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_req
      -- CP-element group 1088: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/$exit
      -- CP-element group 1088: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/$exit
      -- CP-element group 1088: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/$exit
      -- CP-element group 1088: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4139/phi_stmt_4139_sources/type_cast_4142/SplitProtocol/$exit
      -- 
    phi_stmt_4139_req_13665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4139_req_13665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1088), ack => phi_stmt_4139_req_0); -- 
    zeropad3D_cp_element_group_1088: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1088"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1086) & zeropad3D_CP_2152_elements(1087);
      gj_zeropad3D_cp_element_group_1088 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1088), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1089:  transition  input  bypass 
    -- CP-element group 1089: predecessors 
    -- CP-element group 1089: 	602 
    -- CP-element group 1089: successors 
    -- CP-element group 1089: 	1091 
    -- CP-element group 1089:  members (2) 
      -- CP-element group 1089: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Sample/ra
      -- CP-element group 1089: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Sample/$exit
      -- 
    ra_13682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1089_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4148_inst_ack_0, ack => zeropad3D_CP_2152_elements(1089)); -- 
    -- CP-element group 1090:  transition  input  bypass 
    -- CP-element group 1090: predecessors 
    -- CP-element group 1090: 	602 
    -- CP-element group 1090: successors 
    -- CP-element group 1090: 	1091 
    -- CP-element group 1090:  members (2) 
      -- CP-element group 1090: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Update/ca
      -- CP-element group 1090: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/Update/$exit
      -- 
    ca_13687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1090_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4148_inst_ack_1, ack => zeropad3D_CP_2152_elements(1090)); -- 
    -- CP-element group 1091:  join  transition  output  bypass 
    -- CP-element group 1091: predecessors 
    -- CP-element group 1091: 	1089 
    -- CP-element group 1091: 	1090 
    -- CP-element group 1091: successors 
    -- CP-element group 1091: 	1092 
    -- CP-element group 1091:  members (5) 
      -- CP-element group 1091: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/$exit
      -- CP-element group 1091: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_req
      -- CP-element group 1091: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/SplitProtocol/$exit
      -- CP-element group 1091: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/type_cast_4148/$exit
      -- CP-element group 1091: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/phi_stmt_4145/phi_stmt_4145_sources/$exit
      -- 
    phi_stmt_4145_req_13688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4145_req_13688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1091), ack => phi_stmt_4145_req_0); -- 
    zeropad3D_cp_element_group_1091: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1091"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1089) & zeropad3D_CP_2152_elements(1090);
      gj_zeropad3D_cp_element_group_1091 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1091), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1092:  join  transition  bypass 
    -- CP-element group 1092: predecessors 
    -- CP-element group 1092: 	1085 
    -- CP-element group 1092: 	1088 
    -- CP-element group 1092: 	1091 
    -- CP-element group 1092: successors 
    -- CP-element group 1092: 	1093 
    -- CP-element group 1092:  members (1) 
      -- CP-element group 1092: 	 branch_block_stmt_714/ifx_xthen1237_ifx_xend1279_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1092: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1092"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1085) & zeropad3D_CP_2152_elements(1088) & zeropad3D_CP_2152_elements(1091);
      gj_zeropad3D_cp_element_group_1092 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1092), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1093:  merge  fork  transition  place  bypass 
    -- CP-element group 1093: predecessors 
    -- CP-element group 1093: 	1082 
    -- CP-element group 1093: 	1092 
    -- CP-element group 1093: successors 
    -- CP-element group 1093: 	1094 
    -- CP-element group 1093: 	1095 
    -- CP-element group 1093: 	1096 
    -- CP-element group 1093:  members (2) 
      -- CP-element group 1093: 	 branch_block_stmt_714/merge_stmt_4131_PhiReqMerge
      -- CP-element group 1093: 	 branch_block_stmt_714/merge_stmt_4131_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1093) <= OrReduce(zeropad3D_CP_2152_elements(1082) & zeropad3D_CP_2152_elements(1092));
    -- CP-element group 1094:  transition  input  bypass 
    -- CP-element group 1094: predecessors 
    -- CP-element group 1094: 	1093 
    -- CP-element group 1094: successors 
    -- CP-element group 1094: 	1097 
    -- CP-element group 1094:  members (1) 
      -- CP-element group 1094: 	 branch_block_stmt_714/merge_stmt_4131_PhiAck/phi_stmt_4132_ack
      -- 
    phi_stmt_4132_ack_13693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1094_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4132_ack_0, ack => zeropad3D_CP_2152_elements(1094)); -- 
    -- CP-element group 1095:  transition  input  bypass 
    -- CP-element group 1095: predecessors 
    -- CP-element group 1095: 	1093 
    -- CP-element group 1095: successors 
    -- CP-element group 1095: 	1097 
    -- CP-element group 1095:  members (1) 
      -- CP-element group 1095: 	 branch_block_stmt_714/merge_stmt_4131_PhiAck/phi_stmt_4139_ack
      -- 
    phi_stmt_4139_ack_13694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1095_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4139_ack_0, ack => zeropad3D_CP_2152_elements(1095)); -- 
    -- CP-element group 1096:  transition  input  bypass 
    -- CP-element group 1096: predecessors 
    -- CP-element group 1096: 	1093 
    -- CP-element group 1096: successors 
    -- CP-element group 1096: 	1097 
    -- CP-element group 1096:  members (1) 
      -- CP-element group 1096: 	 branch_block_stmt_714/merge_stmt_4131_PhiAck/phi_stmt_4145_ack
      -- 
    phi_stmt_4145_ack_13695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1096_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4145_ack_0, ack => zeropad3D_CP_2152_elements(1096)); -- 
    -- CP-element group 1097:  join  transition  bypass 
    -- CP-element group 1097: predecessors 
    -- CP-element group 1097: 	1094 
    -- CP-element group 1097: 	1095 
    -- CP-element group 1097: 	1096 
    -- CP-element group 1097: successors 
    -- CP-element group 1097: 	6 
    -- CP-element group 1097:  members (1) 
      -- CP-element group 1097: 	 branch_block_stmt_714/merge_stmt_4131_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1097: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1097"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1094) & zeropad3D_CP_2152_elements(1095) & zeropad3D_CP_2152_elements(1096);
      gj_zeropad3D_cp_element_group_1097 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1097), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1098:  transition  input  bypass 
    -- CP-element group 1098: predecessors 
    -- CP-element group 1098: 	7 
    -- CP-element group 1098: successors 
    -- CP-element group 1098: 	1100 
    -- CP-element group 1098:  members (2) 
      -- CP-element group 1098: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Sample/$exit
      -- CP-element group 1098: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Sample/ra
      -- 
    ra_13723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1098_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4303_inst_ack_0, ack => zeropad3D_CP_2152_elements(1098)); -- 
    -- CP-element group 1099:  transition  input  bypass 
    -- CP-element group 1099: predecessors 
    -- CP-element group 1099: 	7 
    -- CP-element group 1099: successors 
    -- CP-element group 1099: 	1100 
    -- CP-element group 1099:  members (2) 
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Update/$exit
      -- CP-element group 1099: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/Update/ca
      -- 
    ca_13728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1099_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4303_inst_ack_1, ack => zeropad3D_CP_2152_elements(1099)); -- 
    -- CP-element group 1100:  join  transition  output  bypass 
    -- CP-element group 1100: predecessors 
    -- CP-element group 1100: 	1098 
    -- CP-element group 1100: 	1099 
    -- CP-element group 1100: successors 
    -- CP-element group 1100: 	1107 
    -- CP-element group 1100:  members (5) 
      -- CP-element group 1100: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_req
      -- CP-element group 1100: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/SplitProtocol/$exit
      -- CP-element group 1100: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4303/$exit
      -- CP-element group 1100: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/$exit
      -- CP-element group 1100: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4297/$exit
      -- 
    phi_stmt_4297_req_13729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4297_req_13729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1100), ack => phi_stmt_4297_req_1); -- 
    zeropad3D_cp_element_group_1100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1098) & zeropad3D_CP_2152_elements(1099);
      gj_zeropad3D_cp_element_group_1100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1101:  transition  input  bypass 
    -- CP-element group 1101: predecessors 
    -- CP-element group 1101: 	7 
    -- CP-element group 1101: successors 
    -- CP-element group 1101: 	1103 
    -- CP-element group 1101:  members (2) 
      -- CP-element group 1101: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Sample/ra
      -- CP-element group 1101: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Sample/$exit
      -- 
    ra_13746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4309_inst_ack_0, ack => zeropad3D_CP_2152_elements(1101)); -- 
    -- CP-element group 1102:  transition  input  bypass 
    -- CP-element group 1102: predecessors 
    -- CP-element group 1102: 	7 
    -- CP-element group 1102: successors 
    -- CP-element group 1102: 	1103 
    -- CP-element group 1102:  members (2) 
      -- CP-element group 1102: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Update/ca
      -- CP-element group 1102: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/Update/$exit
      -- 
    ca_13751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4309_inst_ack_1, ack => zeropad3D_CP_2152_elements(1102)); -- 
    -- CP-element group 1103:  join  transition  output  bypass 
    -- CP-element group 1103: predecessors 
    -- CP-element group 1103: 	1101 
    -- CP-element group 1103: 	1102 
    -- CP-element group 1103: successors 
    -- CP-element group 1103: 	1107 
    -- CP-element group 1103:  members (5) 
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4309/SplitProtocol/$exit
      -- CP-element group 1103: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_req
      -- 
    phi_stmt_4304_req_13752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4304_req_13752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1103), ack => phi_stmt_4304_req_1); -- 
    zeropad3D_cp_element_group_1103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1101) & zeropad3D_CP_2152_elements(1102);
      gj_zeropad3D_cp_element_group_1103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1104:  transition  input  bypass 
    -- CP-element group 1104: predecessors 
    -- CP-element group 1104: 	7 
    -- CP-element group 1104: successors 
    -- CP-element group 1104: 	1106 
    -- CP-element group 1104:  members (2) 
      -- CP-element group 1104: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Sample/$exit
      -- CP-element group 1104: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Sample/ra
      -- 
    ra_13769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4316_inst_ack_0, ack => zeropad3D_CP_2152_elements(1104)); -- 
    -- CP-element group 1105:  transition  input  bypass 
    -- CP-element group 1105: predecessors 
    -- CP-element group 1105: 	7 
    -- CP-element group 1105: successors 
    -- CP-element group 1105: 	1106 
    -- CP-element group 1105:  members (2) 
      -- CP-element group 1105: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Update/$exit
      -- CP-element group 1105: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/Update/ca
      -- 
    ca_13774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4316_inst_ack_1, ack => zeropad3D_CP_2152_elements(1105)); -- 
    -- CP-element group 1106:  join  transition  output  bypass 
    -- CP-element group 1106: predecessors 
    -- CP-element group 1106: 	1104 
    -- CP-element group 1106: 	1105 
    -- CP-element group 1106: successors 
    -- CP-element group 1106: 	1107 
    -- CP-element group 1106:  members (5) 
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/SplitProtocol/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4316/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/$exit
      -- CP-element group 1106: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_req
      -- 
    phi_stmt_4310_req_13775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4310_req_13775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1106), ack => phi_stmt_4310_req_1); -- 
    zeropad3D_cp_element_group_1106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1104) & zeropad3D_CP_2152_elements(1105);
      gj_zeropad3D_cp_element_group_1106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1107:  join  transition  bypass 
    -- CP-element group 1107: predecessors 
    -- CP-element group 1107: 	1100 
    -- CP-element group 1107: 	1103 
    -- CP-element group 1107: 	1106 
    -- CP-element group 1107: successors 
    -- CP-element group 1107: 	1114 
    -- CP-element group 1107:  members (1) 
      -- CP-element group 1107: 	 branch_block_stmt_714/ifx_xend1496_whilex_xbody1341_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1107: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1107"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1100) & zeropad3D_CP_2152_elements(1103) & zeropad3D_CP_2152_elements(1106);
      gj_zeropad3D_cp_element_group_1107 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1108:  transition  output  delay-element  bypass 
    -- CP-element group 1108: predecessors 
    -- CP-element group 1108: 	642 
    -- CP-element group 1108: successors 
    -- CP-element group 1108: 	1113 
    -- CP-element group 1108:  members (4) 
      -- CP-element group 1108: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_req
      -- CP-element group 1108: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/type_cast_4301_konst_delay_trans
      -- CP-element group 1108: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4297/phi_stmt_4297_sources/$exit
      -- CP-element group 1108: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4297/$exit
      -- 
    phi_stmt_4297_req_13786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4297_req_13786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1108), ack => phi_stmt_4297_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1108) is a control-delay.
    cp_element_1108_delay: control_delay_element  generic map(name => " 1108_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(642), ack => zeropad3D_CP_2152_elements(1108), clk => clk, reset =>reset);
    -- CP-element group 1109:  transition  input  bypass 
    -- CP-element group 1109: predecessors 
    -- CP-element group 1109: 	642 
    -- CP-element group 1109: successors 
    -- CP-element group 1109: 	1111 
    -- CP-element group 1109:  members (2) 
      -- CP-element group 1109: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Sample/ra
      -- CP-element group 1109: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Sample/$exit
      -- 
    ra_13803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4307_inst_ack_0, ack => zeropad3D_CP_2152_elements(1109)); -- 
    -- CP-element group 1110:  transition  input  bypass 
    -- CP-element group 1110: predecessors 
    -- CP-element group 1110: 	642 
    -- CP-element group 1110: successors 
    -- CP-element group 1110: 	1111 
    -- CP-element group 1110:  members (2) 
      -- CP-element group 1110: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Update/ca
      -- CP-element group 1110: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/Update/$exit
      -- 
    ca_13808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4307_inst_ack_1, ack => zeropad3D_CP_2152_elements(1110)); -- 
    -- CP-element group 1111:  join  transition  output  bypass 
    -- CP-element group 1111: predecessors 
    -- CP-element group 1111: 	1109 
    -- CP-element group 1111: 	1110 
    -- CP-element group 1111: successors 
    -- CP-element group 1111: 	1113 
    -- CP-element group 1111:  members (5) 
      -- CP-element group 1111: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_req
      -- CP-element group 1111: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/SplitProtocol/$exit
      -- CP-element group 1111: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/type_cast_4307/$exit
      -- CP-element group 1111: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/phi_stmt_4304_sources/$exit
      -- CP-element group 1111: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4304/$exit
      -- 
    phi_stmt_4304_req_13809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4304_req_13809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1111), ack => phi_stmt_4304_req_0); -- 
    zeropad3D_cp_element_group_1111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1109) & zeropad3D_CP_2152_elements(1110);
      gj_zeropad3D_cp_element_group_1111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1112:  transition  output  delay-element  bypass 
    -- CP-element group 1112: predecessors 
    -- CP-element group 1112: 	642 
    -- CP-element group 1112: successors 
    -- CP-element group 1112: 	1113 
    -- CP-element group 1112:  members (4) 
      -- CP-element group 1112: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_req
      -- CP-element group 1112: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/type_cast_4314_konst_delay_trans
      -- CP-element group 1112: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4310/phi_stmt_4310_sources/$exit
      -- CP-element group 1112: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/phi_stmt_4310/$exit
      -- 
    phi_stmt_4310_req_13817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4310_req_13817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1112), ack => phi_stmt_4310_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1112) is a control-delay.
    cp_element_1112_delay: control_delay_element  generic map(name => " 1112_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(642), ack => zeropad3D_CP_2152_elements(1112), clk => clk, reset =>reset);
    -- CP-element group 1113:  join  transition  bypass 
    -- CP-element group 1113: predecessors 
    -- CP-element group 1113: 	1108 
    -- CP-element group 1113: 	1111 
    -- CP-element group 1113: 	1112 
    -- CP-element group 1113: successors 
    -- CP-element group 1113: 	1114 
    -- CP-element group 1113:  members (1) 
      -- CP-element group 1113: 	 branch_block_stmt_714/whilex_xend1280_whilex_xbody1341_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1113: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1113"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1108) & zeropad3D_CP_2152_elements(1111) & zeropad3D_CP_2152_elements(1112);
      gj_zeropad3D_cp_element_group_1113 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1114:  merge  fork  transition  place  bypass 
    -- CP-element group 1114: predecessors 
    -- CP-element group 1114: 	1107 
    -- CP-element group 1114: 	1113 
    -- CP-element group 1114: successors 
    -- CP-element group 1114: 	1115 
    -- CP-element group 1114: 	1116 
    -- CP-element group 1114: 	1117 
    -- CP-element group 1114:  members (2) 
      -- CP-element group 1114: 	 branch_block_stmt_714/merge_stmt_4296_PhiReqMerge
      -- CP-element group 1114: 	 branch_block_stmt_714/merge_stmt_4296_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1114) <= OrReduce(zeropad3D_CP_2152_elements(1107) & zeropad3D_CP_2152_elements(1113));
    -- CP-element group 1115:  transition  input  bypass 
    -- CP-element group 1115: predecessors 
    -- CP-element group 1115: 	1114 
    -- CP-element group 1115: successors 
    -- CP-element group 1115: 	1118 
    -- CP-element group 1115:  members (1) 
      -- CP-element group 1115: 	 branch_block_stmt_714/merge_stmt_4296_PhiAck/phi_stmt_4297_ack
      -- 
    phi_stmt_4297_ack_13822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4297_ack_0, ack => zeropad3D_CP_2152_elements(1115)); -- 
    -- CP-element group 1116:  transition  input  bypass 
    -- CP-element group 1116: predecessors 
    -- CP-element group 1116: 	1114 
    -- CP-element group 1116: successors 
    -- CP-element group 1116: 	1118 
    -- CP-element group 1116:  members (1) 
      -- CP-element group 1116: 	 branch_block_stmt_714/merge_stmt_4296_PhiAck/phi_stmt_4304_ack
      -- 
    phi_stmt_4304_ack_13823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4304_ack_0, ack => zeropad3D_CP_2152_elements(1116)); -- 
    -- CP-element group 1117:  transition  input  bypass 
    -- CP-element group 1117: predecessors 
    -- CP-element group 1117: 	1114 
    -- CP-element group 1117: successors 
    -- CP-element group 1117: 	1118 
    -- CP-element group 1117:  members (1) 
      -- CP-element group 1117: 	 branch_block_stmt_714/merge_stmt_4296_PhiAck/phi_stmt_4310_ack
      -- 
    phi_stmt_4310_ack_13824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4310_ack_0, ack => zeropad3D_CP_2152_elements(1117)); -- 
    -- CP-element group 1118:  join  fork  transition  place  output  bypass 
    -- CP-element group 1118: predecessors 
    -- CP-element group 1118: 	1115 
    -- CP-element group 1118: 	1116 
    -- CP-element group 1118: 	1117 
    -- CP-element group 1118: successors 
    -- CP-element group 1118: 	643 
    -- CP-element group 1118: 	644 
    -- CP-element group 1118:  members (10) 
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329__entry__
      -- CP-element group 1118: 	 branch_block_stmt_714/merge_stmt_4296__exit__
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/$entry
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_sample_start_
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_update_start_
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Sample/$entry
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Sample/rr
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Update/$entry
      -- CP-element group 1118: 	 branch_block_stmt_714/assign_stmt_4322_to_assign_stmt_4329/type_cast_4321_Update/cr
      -- CP-element group 1118: 	 branch_block_stmt_714/merge_stmt_4296_PhiAck/$exit
      -- 
    rr_9617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1118), ack => type_cast_4321_inst_req_0); -- 
    cr_9622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1118), ack => type_cast_4321_inst_req_1); -- 
    zeropad3D_cp_element_group_1118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1115) & zeropad3D_CP_2152_elements(1116) & zeropad3D_CP_2152_elements(1117);
      gj_zeropad3D_cp_element_group_1118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1119:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1119: predecessors 
    -- CP-element group 1119: 	645 
    -- CP-element group 1119: 	652 
    -- CP-element group 1119: 	655 
    -- CP-element group 1119: 	662 
    -- CP-element group 1119: successors 
    -- CP-element group 1119: 	663 
    -- CP-element group 1119: 	664 
    -- CP-element group 1119: 	665 
    -- CP-element group 1119: 	666 
    -- CP-element group 1119: 	669 
    -- CP-element group 1119: 	671 
    -- CP-element group 1119: 	673 
    -- CP-element group 1119: 	675 
    -- CP-element group 1119:  members (33) 
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469__entry__
      -- CP-element group 1119: 	 branch_block_stmt_714/merge_stmt_4413__exit__
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_sample_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_update_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Sample/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Sample/rr
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Update/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4417_Update/cr
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_sample_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_update_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Sample/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Sample/rr
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Update/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4422_Update/cr
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_update_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Update/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/type_cast_4456_Update/cr
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_update_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_update_start
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Update/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/array_obj_ref_4462_final_index_sum_regn_Update/req
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_complete/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/addr_of_4463_complete/req
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_update_start_
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/word_access_complete/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/word_access_complete/word_0/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/assign_stmt_4418_to_assign_stmt_4469/ptr_deref_4466_Update/word_access_complete/word_0/cr
      -- CP-element group 1119: 	 branch_block_stmt_714/merge_stmt_4413_PhiAck/dummy
      -- CP-element group 1119: 	 branch_block_stmt_714/merge_stmt_4413_PhiAck/$exit
      -- CP-element group 1119: 	 branch_block_stmt_714/merge_stmt_4413_PhiAck/$entry
      -- CP-element group 1119: 	 branch_block_stmt_714/merge_stmt_4413_PhiReqMerge
      -- 
    rr_9827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => type_cast_4417_inst_req_0); -- 
    cr_9832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => type_cast_4417_inst_req_1); -- 
    rr_9841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => type_cast_4422_inst_req_0); -- 
    cr_9846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => type_cast_4422_inst_req_1); -- 
    cr_9860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => type_cast_4456_inst_req_1); -- 
    req_9891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => array_obj_ref_4462_index_offset_req_1); -- 
    req_9906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => addr_of_4463_final_reg_req_1); -- 
    cr_9956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1119), ack => ptr_deref_4466_store_0_req_1); -- 
    zeropad3D_CP_2152_elements(1119) <= OrReduce(zeropad3D_CP_2152_elements(645) & zeropad3D_CP_2152_elements(652) & zeropad3D_CP_2152_elements(655) & zeropad3D_CP_2152_elements(662));
    -- CP-element group 1120:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1120: predecessors 
    -- CP-element group 1120: 	676 
    -- CP-element group 1120: 	696 
    -- CP-element group 1120: successors 
    -- CP-element group 1120: 	697 
    -- CP-element group 1120: 	698 
    -- CP-element group 1120:  members (13) 
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596__entry__
      -- CP-element group 1120: 	 branch_block_stmt_714/merge_stmt_4578__exit__
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_sample_start_
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_update_start_
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Sample/rr
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/$entry
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Sample/$entry
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Update/$entry
      -- CP-element group 1120: 	 branch_block_stmt_714/assign_stmt_4583_to_assign_stmt_4596/type_cast_4582_Update/cr
      -- CP-element group 1120: 	 branch_block_stmt_714/merge_stmt_4578_PhiAck/dummy
      -- CP-element group 1120: 	 branch_block_stmt_714/merge_stmt_4578_PhiAck/$exit
      -- CP-element group 1120: 	 branch_block_stmt_714/merge_stmt_4578_PhiAck/$entry
      -- CP-element group 1120: 	 branch_block_stmt_714/merge_stmt_4578_PhiReqMerge
      -- 
    rr_10205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1120), ack => type_cast_4582_inst_req_0); -- 
    cr_10210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1120), ack => type_cast_4582_inst_req_1); -- 
    zeropad3D_CP_2152_elements(1120) <= OrReduce(zeropad3D_CP_2152_elements(676) & zeropad3D_CP_2152_elements(696));
    -- CP-element group 1121:  transition  input  bypass 
    -- CP-element group 1121: predecessors 
    -- CP-element group 1121: 	718 
    -- CP-element group 1121: successors 
    -- CP-element group 1121: 	1123 
    -- CP-element group 1121:  members (2) 
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Sample/ra
      -- CP-element group 1121: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Sample/$exit
      -- 
    ra_13944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4709_inst_ack_0, ack => zeropad3D_CP_2152_elements(1121)); -- 
    -- CP-element group 1122:  transition  input  bypass 
    -- CP-element group 1122: predecessors 
    -- CP-element group 1122: 	718 
    -- CP-element group 1122: successors 
    -- CP-element group 1122: 	1123 
    -- CP-element group 1122:  members (2) 
      -- CP-element group 1122: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Update/ca
      -- CP-element group 1122: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/Update/$exit
      -- 
    ca_13949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4709_inst_ack_1, ack => zeropad3D_CP_2152_elements(1122)); -- 
    -- CP-element group 1123:  join  transition  output  bypass 
    -- CP-element group 1123: predecessors 
    -- CP-element group 1123: 	1121 
    -- CP-element group 1123: 	1122 
    -- CP-element group 1123: successors 
    -- CP-element group 1123: 	1128 
    -- CP-element group 1123:  members (5) 
      -- CP-element group 1123: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_req
      -- CP-element group 1123: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/$exit
      -- CP-element group 1123: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/SplitProtocol/$exit
      -- CP-element group 1123: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4709/$exit
      -- CP-element group 1123: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4704/$exit
      -- 
    phi_stmt_4704_req_13950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4704_req_13950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1123), ack => phi_stmt_4704_req_1); -- 
    zeropad3D_cp_element_group_1123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1121) & zeropad3D_CP_2152_elements(1122);
      gj_zeropad3D_cp_element_group_1123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1124:  transition  input  bypass 
    -- CP-element group 1124: predecessors 
    -- CP-element group 1124: 	718 
    -- CP-element group 1124: successors 
    -- CP-element group 1124: 	1126 
    -- CP-element group 1124:  members (2) 
      -- CP-element group 1124: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Sample/ra
      -- CP-element group 1124: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Sample/$exit
      -- 
    ra_13967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4703_inst_ack_0, ack => zeropad3D_CP_2152_elements(1124)); -- 
    -- CP-element group 1125:  transition  input  bypass 
    -- CP-element group 1125: predecessors 
    -- CP-element group 1125: 	718 
    -- CP-element group 1125: successors 
    -- CP-element group 1125: 	1126 
    -- CP-element group 1125:  members (2) 
      -- CP-element group 1125: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Update/ca
      -- CP-element group 1125: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/Update/$exit
      -- 
    ca_13972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4703_inst_ack_1, ack => zeropad3D_CP_2152_elements(1125)); -- 
    -- CP-element group 1126:  join  transition  output  bypass 
    -- CP-element group 1126: predecessors 
    -- CP-element group 1126: 	1124 
    -- CP-element group 1126: 	1125 
    -- CP-element group 1126: successors 
    -- CP-element group 1126: 	1128 
    -- CP-element group 1126:  members (5) 
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/$exit
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/$exit
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_req
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/SplitProtocol/$exit
      -- CP-element group 1126: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4703/$exit
      -- 
    phi_stmt_4698_req_13973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4698_req_13973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1126), ack => phi_stmt_4698_req_1); -- 
    zeropad3D_cp_element_group_1126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1124) & zeropad3D_CP_2152_elements(1125);
      gj_zeropad3D_cp_element_group_1126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1127:  transition  output  delay-element  bypass 
    -- CP-element group 1127: predecessors 
    -- CP-element group 1127: 	718 
    -- CP-element group 1127: successors 
    -- CP-element group 1127: 	1128 
    -- CP-element group 1127:  members (4) 
      -- CP-element group 1127: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/$exit
      -- CP-element group 1127: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4691/$exit
      -- CP-element group 1127: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_req
      -- CP-element group 1127: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4697_konst_delay_trans
      -- 
    phi_stmt_4691_req_13981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4691_req_13981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1127), ack => phi_stmt_4691_req_1); -- 
    -- Element group zeropad3D_CP_2152_elements(1127) is a control-delay.
    cp_element_1127_delay: control_delay_element  generic map(name => " 1127_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(718), ack => zeropad3D_CP_2152_elements(1127), clk => clk, reset =>reset);
    -- CP-element group 1128:  join  transition  bypass 
    -- CP-element group 1128: predecessors 
    -- CP-element group 1128: 	1123 
    -- CP-element group 1128: 	1126 
    -- CP-element group 1128: 	1127 
    -- CP-element group 1128: successors 
    -- CP-element group 1128: 	1139 
    -- CP-element group 1128:  members (1) 
      -- CP-element group 1128: 	 branch_block_stmt_714/ifx_xelse1460_ifx_xend1496_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1123) & zeropad3D_CP_2152_elements(1126) & zeropad3D_CP_2152_elements(1127);
      gj_zeropad3D_cp_element_group_1128 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1129:  transition  input  bypass 
    -- CP-element group 1129: predecessors 
    -- CP-element group 1129: 	699 
    -- CP-element group 1129: successors 
    -- CP-element group 1129: 	1131 
    -- CP-element group 1129:  members (2) 
      -- CP-element group 1129: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Sample/ra
      -- CP-element group 1129: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Sample/$exit
      -- 
    ra_14001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4707_inst_ack_0, ack => zeropad3D_CP_2152_elements(1129)); -- 
    -- CP-element group 1130:  transition  input  bypass 
    -- CP-element group 1130: predecessors 
    -- CP-element group 1130: 	699 
    -- CP-element group 1130: successors 
    -- CP-element group 1130: 	1131 
    -- CP-element group 1130:  members (2) 
      -- CP-element group 1130: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Update/ca
      -- CP-element group 1130: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/Update/$exit
      -- 
    ca_14006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4707_inst_ack_1, ack => zeropad3D_CP_2152_elements(1130)); -- 
    -- CP-element group 1131:  join  transition  output  bypass 
    -- CP-element group 1131: predecessors 
    -- CP-element group 1131: 	1129 
    -- CP-element group 1131: 	1130 
    -- CP-element group 1131: successors 
    -- CP-element group 1131: 	1138 
    -- CP-element group 1131:  members (5) 
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_req
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/SplitProtocol/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/type_cast_4707/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/phi_stmt_4704_sources/$exit
      -- CP-element group 1131: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4704/$exit
      -- 
    phi_stmt_4704_req_14007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4704_req_14007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1131), ack => phi_stmt_4704_req_0); -- 
    zeropad3D_cp_element_group_1131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1129) & zeropad3D_CP_2152_elements(1130);
      gj_zeropad3D_cp_element_group_1131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1132:  transition  input  bypass 
    -- CP-element group 1132: predecessors 
    -- CP-element group 1132: 	699 
    -- CP-element group 1132: successors 
    -- CP-element group 1132: 	1134 
    -- CP-element group 1132:  members (2) 
      -- CP-element group 1132: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Sample/ra
      -- CP-element group 1132: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Sample/$exit
      -- 
    ra_14024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4701_inst_ack_0, ack => zeropad3D_CP_2152_elements(1132)); -- 
    -- CP-element group 1133:  transition  input  bypass 
    -- CP-element group 1133: predecessors 
    -- CP-element group 1133: 	699 
    -- CP-element group 1133: successors 
    -- CP-element group 1133: 	1134 
    -- CP-element group 1133:  members (2) 
      -- CP-element group 1133: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Update/$exit
      -- CP-element group 1133: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/Update/ca
      -- 
    ca_14029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4701_inst_ack_1, ack => zeropad3D_CP_2152_elements(1133)); -- 
    -- CP-element group 1134:  join  transition  output  bypass 
    -- CP-element group 1134: predecessors 
    -- CP-element group 1134: 	1132 
    -- CP-element group 1134: 	1133 
    -- CP-element group 1134: successors 
    -- CP-element group 1134: 	1138 
    -- CP-element group 1134:  members (5) 
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/SplitProtocol/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_sources/type_cast_4701/$exit
      -- CP-element group 1134: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4698/phi_stmt_4698_req
      -- 
    phi_stmt_4698_req_14030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4698_req_14030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1134), ack => phi_stmt_4698_req_0); -- 
    zeropad3D_cp_element_group_1134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1132) & zeropad3D_CP_2152_elements(1133);
      gj_zeropad3D_cp_element_group_1134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1135:  transition  input  bypass 
    -- CP-element group 1135: predecessors 
    -- CP-element group 1135: 	699 
    -- CP-element group 1135: successors 
    -- CP-element group 1135: 	1137 
    -- CP-element group 1135:  members (2) 
      -- CP-element group 1135: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Sample/$exit
      -- CP-element group 1135: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Sample/ra
      -- 
    ra_14047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4694_inst_ack_0, ack => zeropad3D_CP_2152_elements(1135)); -- 
    -- CP-element group 1136:  transition  input  bypass 
    -- CP-element group 1136: predecessors 
    -- CP-element group 1136: 	699 
    -- CP-element group 1136: successors 
    -- CP-element group 1136: 	1137 
    -- CP-element group 1136:  members (2) 
      -- CP-element group 1136: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Update/$exit
      -- CP-element group 1136: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/Update/ca
      -- 
    ca_14052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4694_inst_ack_1, ack => zeropad3D_CP_2152_elements(1136)); -- 
    -- CP-element group 1137:  join  transition  output  bypass 
    -- CP-element group 1137: predecessors 
    -- CP-element group 1137: 	1135 
    -- CP-element group 1137: 	1136 
    -- CP-element group 1137: successors 
    -- CP-element group 1137: 	1138 
    -- CP-element group 1137:  members (5) 
      -- CP-element group 1137: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/$exit
      -- CP-element group 1137: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/$exit
      -- CP-element group 1137: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/$exit
      -- CP-element group 1137: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_sources/type_cast_4694/SplitProtocol/$exit
      -- CP-element group 1137: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/phi_stmt_4691/phi_stmt_4691_req
      -- 
    phi_stmt_4691_req_14053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4691_req_14053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1137), ack => phi_stmt_4691_req_0); -- 
    zeropad3D_cp_element_group_1137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1135) & zeropad3D_CP_2152_elements(1136);
      gj_zeropad3D_cp_element_group_1137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1138:  join  transition  bypass 
    -- CP-element group 1138: predecessors 
    -- CP-element group 1138: 	1131 
    -- CP-element group 1138: 	1134 
    -- CP-element group 1138: 	1137 
    -- CP-element group 1138: successors 
    -- CP-element group 1138: 	1139 
    -- CP-element group 1138:  members (1) 
      -- CP-element group 1138: 	 branch_block_stmt_714/ifx_xthen1455_ifx_xend1496_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1138: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1138"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1131) & zeropad3D_CP_2152_elements(1134) & zeropad3D_CP_2152_elements(1137);
      gj_zeropad3D_cp_element_group_1138 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1139:  merge  fork  transition  place  bypass 
    -- CP-element group 1139: predecessors 
    -- CP-element group 1139: 	1128 
    -- CP-element group 1139: 	1138 
    -- CP-element group 1139: successors 
    -- CP-element group 1139: 	1140 
    -- CP-element group 1139: 	1141 
    -- CP-element group 1139: 	1142 
    -- CP-element group 1139:  members (2) 
      -- CP-element group 1139: 	 branch_block_stmt_714/merge_stmt_4690_PhiReqMerge
      -- CP-element group 1139: 	 branch_block_stmt_714/merge_stmt_4690_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1139) <= OrReduce(zeropad3D_CP_2152_elements(1128) & zeropad3D_CP_2152_elements(1138));
    -- CP-element group 1140:  transition  input  bypass 
    -- CP-element group 1140: predecessors 
    -- CP-element group 1140: 	1139 
    -- CP-element group 1140: successors 
    -- CP-element group 1140: 	1143 
    -- CP-element group 1140:  members (1) 
      -- CP-element group 1140: 	 branch_block_stmt_714/merge_stmt_4690_PhiAck/phi_stmt_4691_ack
      -- 
    phi_stmt_4691_ack_14058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4691_ack_0, ack => zeropad3D_CP_2152_elements(1140)); -- 
    -- CP-element group 1141:  transition  input  bypass 
    -- CP-element group 1141: predecessors 
    -- CP-element group 1141: 	1139 
    -- CP-element group 1141: successors 
    -- CP-element group 1141: 	1143 
    -- CP-element group 1141:  members (1) 
      -- CP-element group 1141: 	 branch_block_stmt_714/merge_stmt_4690_PhiAck/phi_stmt_4698_ack
      -- 
    phi_stmt_4698_ack_14059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4698_ack_0, ack => zeropad3D_CP_2152_elements(1141)); -- 
    -- CP-element group 1142:  transition  input  bypass 
    -- CP-element group 1142: predecessors 
    -- CP-element group 1142: 	1139 
    -- CP-element group 1142: successors 
    -- CP-element group 1142: 	1143 
    -- CP-element group 1142:  members (1) 
      -- CP-element group 1142: 	 branch_block_stmt_714/merge_stmt_4690_PhiAck/phi_stmt_4704_ack
      -- 
    phi_stmt_4704_ack_14060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4704_ack_0, ack => zeropad3D_CP_2152_elements(1142)); -- 
    -- CP-element group 1143:  join  transition  bypass 
    -- CP-element group 1143: predecessors 
    -- CP-element group 1143: 	1140 
    -- CP-element group 1143: 	1141 
    -- CP-element group 1143: 	1142 
    -- CP-element group 1143: successors 
    -- CP-element group 1143: 	7 
    -- CP-element group 1143:  members (1) 
      -- CP-element group 1143: 	 branch_block_stmt_714/merge_stmt_4690_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1143: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1143"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1140) & zeropad3D_CP_2152_elements(1141) & zeropad3D_CP_2152_elements(1142);
      gj_zeropad3D_cp_element_group_1143 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1144:  transition  input  bypass 
    -- CP-element group 1144: predecessors 
    -- CP-element group 1144: 	8 
    -- CP-element group 1144: successors 
    -- CP-element group 1144: 	1146 
    -- CP-element group 1144:  members (2) 
      -- CP-element group 1144: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Sample/$exit
      -- CP-element group 1144: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Sample/ra
      -- 
    ra_14088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4884_inst_ack_0, ack => zeropad3D_CP_2152_elements(1144)); -- 
    -- CP-element group 1145:  transition  input  bypass 
    -- CP-element group 1145: predecessors 
    -- CP-element group 1145: 	8 
    -- CP-element group 1145: successors 
    -- CP-element group 1145: 	1146 
    -- CP-element group 1145:  members (2) 
      -- CP-element group 1145: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Update/$exit
      -- CP-element group 1145: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/Update/ca
      -- 
    ca_14093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4884_inst_ack_1, ack => zeropad3D_CP_2152_elements(1145)); -- 
    -- CP-element group 1146:  join  transition  output  bypass 
    -- CP-element group 1146: predecessors 
    -- CP-element group 1146: 	1144 
    -- CP-element group 1146: 	1145 
    -- CP-element group 1146: successors 
    -- CP-element group 1146: 	1153 
    -- CP-element group 1146:  members (5) 
      -- CP-element group 1146: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/$exit
      -- CP-element group 1146: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/$exit
      -- CP-element group 1146: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/$exit
      -- CP-element group 1146: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4884/SplitProtocol/$exit
      -- CP-element group 1146: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_req
      -- 
    phi_stmt_4879_req_14094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4879_req_14094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1146), ack => phi_stmt_4879_req_1); -- 
    zeropad3D_cp_element_group_1146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1144) & zeropad3D_CP_2152_elements(1145);
      gj_zeropad3D_cp_element_group_1146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1147:  transition  input  bypass 
    -- CP-element group 1147: predecessors 
    -- CP-element group 1147: 	8 
    -- CP-element group 1147: successors 
    -- CP-element group 1147: 	1149 
    -- CP-element group 1147:  members (2) 
      -- CP-element group 1147: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Sample/$exit
      -- CP-element group 1147: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Sample/ra
      -- 
    ra_14111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4876_inst_ack_0, ack => zeropad3D_CP_2152_elements(1147)); -- 
    -- CP-element group 1148:  transition  input  bypass 
    -- CP-element group 1148: predecessors 
    -- CP-element group 1148: 	8 
    -- CP-element group 1148: successors 
    -- CP-element group 1148: 	1149 
    -- CP-element group 1148:  members (2) 
      -- CP-element group 1148: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Update/$exit
      -- CP-element group 1148: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/Update/ca
      -- 
    ca_14116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4876_inst_ack_1, ack => zeropad3D_CP_2152_elements(1148)); -- 
    -- CP-element group 1149:  join  transition  output  bypass 
    -- CP-element group 1149: predecessors 
    -- CP-element group 1149: 	1147 
    -- CP-element group 1149: 	1148 
    -- CP-element group 1149: successors 
    -- CP-element group 1149: 	1153 
    -- CP-element group 1149:  members (5) 
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/$exit
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/$exit
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/$exit
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4876/SplitProtocol/$exit
      -- CP-element group 1149: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_req
      -- 
    phi_stmt_4873_req_14117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4873_req_14117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1149), ack => phi_stmt_4873_req_0); -- 
    zeropad3D_cp_element_group_1149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1147) & zeropad3D_CP_2152_elements(1148);
      gj_zeropad3D_cp_element_group_1149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1150:  transition  input  bypass 
    -- CP-element group 1150: predecessors 
    -- CP-element group 1150: 	8 
    -- CP-element group 1150: successors 
    -- CP-element group 1150: 	1152 
    -- CP-element group 1150:  members (2) 
      -- CP-element group 1150: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Sample/$exit
      -- CP-element group 1150: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Sample/ra
      -- 
    ra_14134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4872_inst_ack_0, ack => zeropad3D_CP_2152_elements(1150)); -- 
    -- CP-element group 1151:  transition  input  bypass 
    -- CP-element group 1151: predecessors 
    -- CP-element group 1151: 	8 
    -- CP-element group 1151: successors 
    -- CP-element group 1151: 	1152 
    -- CP-element group 1151:  members (2) 
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Update/$exit
      -- CP-element group 1151: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/Update/ca
      -- 
    ca_14139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4872_inst_ack_1, ack => zeropad3D_CP_2152_elements(1151)); -- 
    -- CP-element group 1152:  join  transition  output  bypass 
    -- CP-element group 1152: predecessors 
    -- CP-element group 1152: 	1150 
    -- CP-element group 1152: 	1151 
    -- CP-element group 1152: successors 
    -- CP-element group 1152: 	1153 
    -- CP-element group 1152:  members (5) 
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/$exit
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/$exit
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/$exit
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4872/SplitProtocol/$exit
      -- CP-element group 1152: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_req
      -- 
    phi_stmt_4866_req_14140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4866_req_14140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1152), ack => phi_stmt_4866_req_1); -- 
    zeropad3D_cp_element_group_1152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1150) & zeropad3D_CP_2152_elements(1151);
      gj_zeropad3D_cp_element_group_1152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1153:  join  transition  bypass 
    -- CP-element group 1153: predecessors 
    -- CP-element group 1153: 	1146 
    -- CP-element group 1153: 	1149 
    -- CP-element group 1153: 	1152 
    -- CP-element group 1153: successors 
    -- CP-element group 1153: 	1162 
    -- CP-element group 1153:  members (1) 
      -- CP-element group 1153: 	 branch_block_stmt_714/ifx_xend1715_whilex_xbody1562_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1153: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1153"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1146) & zeropad3D_CP_2152_elements(1149) & zeropad3D_CP_2152_elements(1152);
      gj_zeropad3D_cp_element_group_1153 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1154:  transition  input  bypass 
    -- CP-element group 1154: predecessors 
    -- CP-element group 1154: 	741 
    -- CP-element group 1154: successors 
    -- CP-element group 1154: 	1156 
    -- CP-element group 1154:  members (2) 
      -- CP-element group 1154: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Sample/$exit
      -- CP-element group 1154: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Sample/ra
      -- 
    ra_14160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4882_inst_ack_0, ack => zeropad3D_CP_2152_elements(1154)); -- 
    -- CP-element group 1155:  transition  input  bypass 
    -- CP-element group 1155: predecessors 
    -- CP-element group 1155: 	741 
    -- CP-element group 1155: successors 
    -- CP-element group 1155: 	1156 
    -- CP-element group 1155:  members (2) 
      -- CP-element group 1155: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Update/$exit
      -- CP-element group 1155: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/Update/ca
      -- 
    ca_14165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4882_inst_ack_1, ack => zeropad3D_CP_2152_elements(1155)); -- 
    -- CP-element group 1156:  join  transition  output  bypass 
    -- CP-element group 1156: predecessors 
    -- CP-element group 1156: 	1154 
    -- CP-element group 1156: 	1155 
    -- CP-element group 1156: successors 
    -- CP-element group 1156: 	1161 
    -- CP-element group 1156:  members (5) 
      -- CP-element group 1156: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/$exit
      -- CP-element group 1156: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/$exit
      -- CP-element group 1156: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/$exit
      -- CP-element group 1156: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_sources/type_cast_4882/SplitProtocol/$exit
      -- CP-element group 1156: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4879/phi_stmt_4879_req
      -- 
    phi_stmt_4879_req_14166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4879_req_14166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1156), ack => phi_stmt_4879_req_0); -- 
    zeropad3D_cp_element_group_1156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1154) & zeropad3D_CP_2152_elements(1155);
      gj_zeropad3D_cp_element_group_1156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1157:  transition  input  bypass 
    -- CP-element group 1157: predecessors 
    -- CP-element group 1157: 	741 
    -- CP-element group 1157: successors 
    -- CP-element group 1157: 	1159 
    -- CP-element group 1157:  members (2) 
      -- CP-element group 1157: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Sample/$exit
      -- CP-element group 1157: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Sample/ra
      -- 
    ra_14183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4878_inst_ack_0, ack => zeropad3D_CP_2152_elements(1157)); -- 
    -- CP-element group 1158:  transition  input  bypass 
    -- CP-element group 1158: predecessors 
    -- CP-element group 1158: 	741 
    -- CP-element group 1158: successors 
    -- CP-element group 1158: 	1159 
    -- CP-element group 1158:  members (2) 
      -- CP-element group 1158: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Update/$exit
      -- CP-element group 1158: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/Update/ca
      -- 
    ca_14188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_4878_inst_ack_1, ack => zeropad3D_CP_2152_elements(1158)); -- 
    -- CP-element group 1159:  join  transition  output  bypass 
    -- CP-element group 1159: predecessors 
    -- CP-element group 1159: 	1157 
    -- CP-element group 1159: 	1158 
    -- CP-element group 1159: successors 
    -- CP-element group 1159: 	1161 
    -- CP-element group 1159:  members (5) 
      -- CP-element group 1159: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_sources/type_cast_4878/SplitProtocol/$exit
      -- CP-element group 1159: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4873/phi_stmt_4873_req
      -- 
    phi_stmt_4873_req_14189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4873_req_14189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1159), ack => phi_stmt_4873_req_1); -- 
    zeropad3D_cp_element_group_1159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1157) & zeropad3D_CP_2152_elements(1158);
      gj_zeropad3D_cp_element_group_1159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1160:  transition  output  delay-element  bypass 
    -- CP-element group 1160: predecessors 
    -- CP-element group 1160: 	741 
    -- CP-element group 1160: successors 
    -- CP-element group 1160: 	1161 
    -- CP-element group 1160:  members (4) 
      -- CP-element group 1160: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4866/$exit
      -- CP-element group 1160: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/$exit
      -- CP-element group 1160: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_sources/type_cast_4870_konst_delay_trans
      -- CP-element group 1160: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/phi_stmt_4866/phi_stmt_4866_req
      -- 
    phi_stmt_4866_req_14197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4866_req_14197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1160), ack => phi_stmt_4866_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1160) is a control-delay.
    cp_element_1160_delay: control_delay_element  generic map(name => " 1160_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(741), ack => zeropad3D_CP_2152_elements(1160), clk => clk, reset =>reset);
    -- CP-element group 1161:  join  transition  bypass 
    -- CP-element group 1161: predecessors 
    -- CP-element group 1161: 	1156 
    -- CP-element group 1161: 	1159 
    -- CP-element group 1161: 	1160 
    -- CP-element group 1161: successors 
    -- CP-element group 1161: 	1162 
    -- CP-element group 1161:  members (1) 
      -- CP-element group 1161: 	 branch_block_stmt_714/whilex_xend1497_whilex_xbody1562_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1161: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1161"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1156) & zeropad3D_CP_2152_elements(1159) & zeropad3D_CP_2152_elements(1160);
      gj_zeropad3D_cp_element_group_1161 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1162:  merge  fork  transition  place  bypass 
    -- CP-element group 1162: predecessors 
    -- CP-element group 1162: 	1153 
    -- CP-element group 1162: 	1161 
    -- CP-element group 1162: successors 
    -- CP-element group 1162: 	1163 
    -- CP-element group 1162: 	1164 
    -- CP-element group 1162: 	1165 
    -- CP-element group 1162:  members (2) 
      -- CP-element group 1162: 	 branch_block_stmt_714/merge_stmt_4865_PhiReqMerge
      -- CP-element group 1162: 	 branch_block_stmt_714/merge_stmt_4865_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1162) <= OrReduce(zeropad3D_CP_2152_elements(1153) & zeropad3D_CP_2152_elements(1161));
    -- CP-element group 1163:  transition  input  bypass 
    -- CP-element group 1163: predecessors 
    -- CP-element group 1163: 	1162 
    -- CP-element group 1163: successors 
    -- CP-element group 1163: 	1166 
    -- CP-element group 1163:  members (1) 
      -- CP-element group 1163: 	 branch_block_stmt_714/merge_stmt_4865_PhiAck/phi_stmt_4866_ack
      -- 
    phi_stmt_4866_ack_14202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4866_ack_0, ack => zeropad3D_CP_2152_elements(1163)); -- 
    -- CP-element group 1164:  transition  input  bypass 
    -- CP-element group 1164: predecessors 
    -- CP-element group 1164: 	1162 
    -- CP-element group 1164: successors 
    -- CP-element group 1164: 	1166 
    -- CP-element group 1164:  members (1) 
      -- CP-element group 1164: 	 branch_block_stmt_714/merge_stmt_4865_PhiAck/phi_stmt_4873_ack
      -- 
    phi_stmt_4873_ack_14203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4873_ack_0, ack => zeropad3D_CP_2152_elements(1164)); -- 
    -- CP-element group 1165:  transition  input  bypass 
    -- CP-element group 1165: predecessors 
    -- CP-element group 1165: 	1162 
    -- CP-element group 1165: successors 
    -- CP-element group 1165: 	1166 
    -- CP-element group 1165:  members (1) 
      -- CP-element group 1165: 	 branch_block_stmt_714/merge_stmt_4865_PhiAck/phi_stmt_4879_ack
      -- 
    phi_stmt_4879_ack_14204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4879_ack_0, ack => zeropad3D_CP_2152_elements(1165)); -- 
    -- CP-element group 1166:  join  fork  transition  place  output  bypass 
    -- CP-element group 1166: predecessors 
    -- CP-element group 1166: 	1163 
    -- CP-element group 1166: 	1164 
    -- CP-element group 1166: 	1165 
    -- CP-element group 1166: successors 
    -- CP-element group 1166: 	742 
    -- CP-element group 1166: 	743 
    -- CP-element group 1166:  members (10) 
      -- CP-element group 1166: 	 branch_block_stmt_714/merge_stmt_4865__exit__
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897__entry__
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/$entry
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_sample_start_
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_update_start_
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Sample/$entry
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Sample/rr
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Update/$entry
      -- CP-element group 1166: 	 branch_block_stmt_714/assign_stmt_4890_to_assign_stmt_4897/type_cast_4889_Update/cr
      -- CP-element group 1166: 	 branch_block_stmt_714/merge_stmt_4865_PhiAck/$exit
      -- 
    rr_10707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1166), ack => type_cast_4889_inst_req_0); -- 
    cr_10712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1166), ack => type_cast_4889_inst_req_1); -- 
    zeropad3D_cp_element_group_1166: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1166"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1163) & zeropad3D_CP_2152_elements(1164) & zeropad3D_CP_2152_elements(1165);
      gj_zeropad3D_cp_element_group_1166 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1167:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1167: predecessors 
    -- CP-element group 1167: 	744 
    -- CP-element group 1167: 	751 
    -- CP-element group 1167: 	754 
    -- CP-element group 1167: 	761 
    -- CP-element group 1167: successors 
    -- CP-element group 1167: 	762 
    -- CP-element group 1167: 	763 
    -- CP-element group 1167: 	764 
    -- CP-element group 1167: 	765 
    -- CP-element group 1167: 	768 
    -- CP-element group 1167: 	770 
    -- CP-element group 1167: 	772 
    -- CP-element group 1167: 	774 
    -- CP-element group 1167:  members (33) 
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4975__exit__
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031__entry__
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_update_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_update_start
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Update/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/array_obj_ref_5024_final_index_sum_regn_Update/req
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_sample_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_update_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Update/cr
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_Update/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_update_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_5018_update_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Update/cr
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_complete/req
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Update/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/word_access_complete/word_0/cr
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Sample/rr
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_Sample/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/word_access_complete/word_0/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/word_access_complete/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/ptr_deref_5028_Update/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_update_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4984_sample_start_
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/addr_of_5025_complete/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Update/cr
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Update/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Sample/rr
      -- CP-element group 1167: 	 branch_block_stmt_714/assign_stmt_4980_to_assign_stmt_5031/type_cast_4979_Sample/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4975_PhiReqMerge
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4975_PhiAck/$entry
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4975_PhiAck/$exit
      -- CP-element group 1167: 	 branch_block_stmt_714/merge_stmt_4975_PhiAck/dummy
      -- 
    req_10981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => array_obj_ref_5024_index_offset_req_1); -- 
    cr_10950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => type_cast_5018_inst_req_1); -- 
    cr_10936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => type_cast_4984_inst_req_1); -- 
    req_10996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => addr_of_5025_final_reg_req_1); -- 
    cr_11046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => ptr_deref_5028_store_0_req_1); -- 
    rr_10931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => type_cast_4984_inst_req_0); -- 
    cr_10922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => type_cast_4979_inst_req_1); -- 
    rr_10917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1167), ack => type_cast_4979_inst_req_0); -- 
    zeropad3D_CP_2152_elements(1167) <= OrReduce(zeropad3D_CP_2152_elements(744) & zeropad3D_CP_2152_elements(751) & zeropad3D_CP_2152_elements(754) & zeropad3D_CP_2152_elements(761));
    -- CP-element group 1168:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1168: predecessors 
    -- CP-element group 1168: 	775 
    -- CP-element group 1168: 	795 
    -- CP-element group 1168: successors 
    -- CP-element group 1168: 	796 
    -- CP-element group 1168: 	797 
    -- CP-element group 1168:  members (13) 
      -- CP-element group 1168: 	 branch_block_stmt_714/merge_stmt_5140__exit__
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158__entry__
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/$entry
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Update/cr
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Update/$entry
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Sample/rr
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_Sample/$entry
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_update_start_
      -- CP-element group 1168: 	 branch_block_stmt_714/assign_stmt_5145_to_assign_stmt_5158/type_cast_5144_sample_start_
      -- CP-element group 1168: 	 branch_block_stmt_714/merge_stmt_5140_PhiReqMerge
      -- CP-element group 1168: 	 branch_block_stmt_714/merge_stmt_5140_PhiAck/$entry
      -- CP-element group 1168: 	 branch_block_stmt_714/merge_stmt_5140_PhiAck/$exit
      -- CP-element group 1168: 	 branch_block_stmt_714/merge_stmt_5140_PhiAck/dummy
      -- 
    cr_11300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_11300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1168), ack => type_cast_5144_inst_req_1); -- 
    rr_11295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_11295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1168), ack => type_cast_5144_inst_req_0); -- 
    zeropad3D_CP_2152_elements(1168) <= OrReduce(zeropad3D_CP_2152_elements(775) & zeropad3D_CP_2152_elements(795));
    -- CP-element group 1169:  transition  output  delay-element  bypass 
    -- CP-element group 1169: predecessors 
    -- CP-element group 1169: 	817 
    -- CP-element group 1169: successors 
    -- CP-element group 1169: 	1176 
    -- CP-element group 1169:  members (4) 
      -- CP-element group 1169: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5246/$exit
      -- CP-element group 1169: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/$exit
      -- CP-element group 1169: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5250_konst_delay_trans
      -- CP-element group 1169: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_req
      -- 
    phi_stmt_5246_req_14315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5246_req_14315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1169), ack => phi_stmt_5246_req_0); -- 
    -- Element group zeropad3D_CP_2152_elements(1169) is a control-delay.
    cp_element_1169_delay: control_delay_element  generic map(name => " 1169_delay", delay_value => 1)  port map(req => zeropad3D_CP_2152_elements(817), ack => zeropad3D_CP_2152_elements(1169), clk => clk, reset =>reset);
    -- CP-element group 1170:  transition  input  bypass 
    -- CP-element group 1170: predecessors 
    -- CP-element group 1170: 	817 
    -- CP-element group 1170: successors 
    -- CP-element group 1170: 	1172 
    -- CP-element group 1170:  members (2) 
      -- CP-element group 1170: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Sample/$exit
      -- CP-element group 1170: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Sample/ra
      -- 
    ra_14332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5258_inst_ack_0, ack => zeropad3D_CP_2152_elements(1170)); -- 
    -- CP-element group 1171:  transition  input  bypass 
    -- CP-element group 1171: predecessors 
    -- CP-element group 1171: 	817 
    -- CP-element group 1171: successors 
    -- CP-element group 1171: 	1172 
    -- CP-element group 1171:  members (2) 
      -- CP-element group 1171: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Update/$exit
      -- CP-element group 1171: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/Update/ca
      -- 
    ca_14337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5258_inst_ack_1, ack => zeropad3D_CP_2152_elements(1171)); -- 
    -- CP-element group 1172:  join  transition  output  bypass 
    -- CP-element group 1172: predecessors 
    -- CP-element group 1172: 	1170 
    -- CP-element group 1172: 	1171 
    -- CP-element group 1172: successors 
    -- CP-element group 1172: 	1176 
    -- CP-element group 1172:  members (5) 
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/$exit
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/$exit
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/$exit
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5258/SplitProtocol/$exit
      -- CP-element group 1172: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_req
      -- 
    phi_stmt_5253_req_14338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5253_req_14338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1172), ack => phi_stmt_5253_req_1); -- 
    zeropad3D_cp_element_group_1172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1170) & zeropad3D_CP_2152_elements(1171);
      gj_zeropad3D_cp_element_group_1172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1173:  transition  input  bypass 
    -- CP-element group 1173: predecessors 
    -- CP-element group 1173: 	817 
    -- CP-element group 1173: successors 
    -- CP-element group 1173: 	1175 
    -- CP-element group 1173:  members (2) 
      -- CP-element group 1173: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Sample/$exit
      -- CP-element group 1173: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Sample/ra
      -- 
    ra_14355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5264_inst_ack_0, ack => zeropad3D_CP_2152_elements(1173)); -- 
    -- CP-element group 1174:  transition  input  bypass 
    -- CP-element group 1174: predecessors 
    -- CP-element group 1174: 	817 
    -- CP-element group 1174: successors 
    -- CP-element group 1174: 	1175 
    -- CP-element group 1174:  members (2) 
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Update/$exit
      -- CP-element group 1174: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/Update/ca
      -- 
    ca_14360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5264_inst_ack_1, ack => zeropad3D_CP_2152_elements(1174)); -- 
    -- CP-element group 1175:  join  transition  output  bypass 
    -- CP-element group 1175: predecessors 
    -- CP-element group 1175: 	1173 
    -- CP-element group 1175: 	1174 
    -- CP-element group 1175: successors 
    -- CP-element group 1175: 	1176 
    -- CP-element group 1175:  members (5) 
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/$exit
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/$exit
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/$exit
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5264/SplitProtocol/$exit
      -- CP-element group 1175: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_req
      -- 
    phi_stmt_5259_req_14361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5259_req_14361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1175), ack => phi_stmt_5259_req_1); -- 
    zeropad3D_cp_element_group_1175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1173) & zeropad3D_CP_2152_elements(1174);
      gj_zeropad3D_cp_element_group_1175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1176:  join  transition  bypass 
    -- CP-element group 1176: predecessors 
    -- CP-element group 1176: 	1169 
    -- CP-element group 1176: 	1172 
    -- CP-element group 1176: 	1175 
    -- CP-element group 1176: successors 
    -- CP-element group 1176: 	1187 
    -- CP-element group 1176:  members (1) 
      -- CP-element group 1176: 	 branch_block_stmt_714/ifx_xelse1680_ifx_xend1715_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1176: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1176"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1169) & zeropad3D_CP_2152_elements(1172) & zeropad3D_CP_2152_elements(1175);
      gj_zeropad3D_cp_element_group_1176 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1177:  transition  input  bypass 
    -- CP-element group 1177: predecessors 
    -- CP-element group 1177: 	798 
    -- CP-element group 1177: successors 
    -- CP-element group 1177: 	1179 
    -- CP-element group 1177:  members (2) 
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Sample/$exit
      -- CP-element group 1177: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Sample/ra
      -- 
    ra_14381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5252_inst_ack_0, ack => zeropad3D_CP_2152_elements(1177)); -- 
    -- CP-element group 1178:  transition  input  bypass 
    -- CP-element group 1178: predecessors 
    -- CP-element group 1178: 	798 
    -- CP-element group 1178: successors 
    -- CP-element group 1178: 	1179 
    -- CP-element group 1178:  members (2) 
      -- CP-element group 1178: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Update/$exit
      -- CP-element group 1178: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/Update/ca
      -- 
    ca_14386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5252_inst_ack_1, ack => zeropad3D_CP_2152_elements(1178)); -- 
    -- CP-element group 1179:  join  transition  output  bypass 
    -- CP-element group 1179: predecessors 
    -- CP-element group 1179: 	1177 
    -- CP-element group 1179: 	1178 
    -- CP-element group 1179: successors 
    -- CP-element group 1179: 	1186 
    -- CP-element group 1179:  members (5) 
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/$exit
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/$exit
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/$exit
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_sources/type_cast_5252/SplitProtocol/$exit
      -- CP-element group 1179: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5246/phi_stmt_5246_req
      -- 
    phi_stmt_5246_req_14387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5246_req_14387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1179), ack => phi_stmt_5246_req_1); -- 
    zeropad3D_cp_element_group_1179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1177) & zeropad3D_CP_2152_elements(1178);
      gj_zeropad3D_cp_element_group_1179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1180:  transition  input  bypass 
    -- CP-element group 1180: predecessors 
    -- CP-element group 1180: 	798 
    -- CP-element group 1180: successors 
    -- CP-element group 1180: 	1182 
    -- CP-element group 1180:  members (2) 
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Sample/$exit
      -- CP-element group 1180: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Sample/ra
      -- 
    ra_14404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5256_inst_ack_0, ack => zeropad3D_CP_2152_elements(1180)); -- 
    -- CP-element group 1181:  transition  input  bypass 
    -- CP-element group 1181: predecessors 
    -- CP-element group 1181: 	798 
    -- CP-element group 1181: successors 
    -- CP-element group 1181: 	1182 
    -- CP-element group 1181:  members (2) 
      -- CP-element group 1181: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Update/$exit
      -- CP-element group 1181: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/Update/ca
      -- 
    ca_14409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5256_inst_ack_1, ack => zeropad3D_CP_2152_elements(1181)); -- 
    -- CP-element group 1182:  join  transition  output  bypass 
    -- CP-element group 1182: predecessors 
    -- CP-element group 1182: 	1180 
    -- CP-element group 1182: 	1181 
    -- CP-element group 1182: successors 
    -- CP-element group 1182: 	1186 
    -- CP-element group 1182:  members (5) 
      -- CP-element group 1182: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/$exit
      -- CP-element group 1182: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/$exit
      -- CP-element group 1182: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/$exit
      -- CP-element group 1182: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_sources/type_cast_5256/SplitProtocol/$exit
      -- CP-element group 1182: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5253/phi_stmt_5253_req
      -- 
    phi_stmt_5253_req_14410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5253_req_14410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1182), ack => phi_stmt_5253_req_0); -- 
    zeropad3D_cp_element_group_1182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1180) & zeropad3D_CP_2152_elements(1181);
      gj_zeropad3D_cp_element_group_1182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1183:  transition  input  bypass 
    -- CP-element group 1183: predecessors 
    -- CP-element group 1183: 	798 
    -- CP-element group 1183: successors 
    -- CP-element group 1183: 	1185 
    -- CP-element group 1183:  members (2) 
      -- CP-element group 1183: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Sample/$exit
      -- CP-element group 1183: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Sample/ra
      -- 
    ra_14427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5262_inst_ack_0, ack => zeropad3D_CP_2152_elements(1183)); -- 
    -- CP-element group 1184:  transition  input  bypass 
    -- CP-element group 1184: predecessors 
    -- CP-element group 1184: 	798 
    -- CP-element group 1184: successors 
    -- CP-element group 1184: 	1185 
    -- CP-element group 1184:  members (2) 
      -- CP-element group 1184: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Update/$exit
      -- CP-element group 1184: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/Update/ca
      -- 
    ca_14432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_5262_inst_ack_1, ack => zeropad3D_CP_2152_elements(1184)); -- 
    -- CP-element group 1185:  join  transition  output  bypass 
    -- CP-element group 1185: predecessors 
    -- CP-element group 1185: 	1183 
    -- CP-element group 1185: 	1184 
    -- CP-element group 1185: successors 
    -- CP-element group 1185: 	1186 
    -- CP-element group 1185:  members (5) 
      -- CP-element group 1185: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_sources/type_cast_5262/SplitProtocol/$exit
      -- CP-element group 1185: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/phi_stmt_5259/phi_stmt_5259_req
      -- 
    phi_stmt_5259_req_14433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_5259_req_14433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_2152_elements(1185), ack => phi_stmt_5259_req_0); -- 
    zeropad3D_cp_element_group_1185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1183) & zeropad3D_CP_2152_elements(1184);
      gj_zeropad3D_cp_element_group_1185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1186:  join  transition  bypass 
    -- CP-element group 1186: predecessors 
    -- CP-element group 1186: 	1179 
    -- CP-element group 1186: 	1182 
    -- CP-element group 1186: 	1185 
    -- CP-element group 1186: successors 
    -- CP-element group 1186: 	1187 
    -- CP-element group 1186:  members (1) 
      -- CP-element group 1186: 	 branch_block_stmt_714/ifx_xthen1675_ifx_xend1715_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_1186: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1186"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1179) & zeropad3D_CP_2152_elements(1182) & zeropad3D_CP_2152_elements(1185);
      gj_zeropad3D_cp_element_group_1186 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 1187:  merge  fork  transition  place  bypass 
    -- CP-element group 1187: predecessors 
    -- CP-element group 1187: 	1176 
    -- CP-element group 1187: 	1186 
    -- CP-element group 1187: successors 
    -- CP-element group 1187: 	1188 
    -- CP-element group 1187: 	1189 
    -- CP-element group 1187: 	1190 
    -- CP-element group 1187:  members (2) 
      -- CP-element group 1187: 	 branch_block_stmt_714/merge_stmt_5245_PhiReqMerge
      -- CP-element group 1187: 	 branch_block_stmt_714/merge_stmt_5245_PhiAck/$entry
      -- 
    zeropad3D_CP_2152_elements(1187) <= OrReduce(zeropad3D_CP_2152_elements(1176) & zeropad3D_CP_2152_elements(1186));
    -- CP-element group 1188:  transition  input  bypass 
    -- CP-element group 1188: predecessors 
    -- CP-element group 1188: 	1187 
    -- CP-element group 1188: successors 
    -- CP-element group 1188: 	1191 
    -- CP-element group 1188:  members (1) 
      -- CP-element group 1188: 	 branch_block_stmt_714/merge_stmt_5245_PhiAck/phi_stmt_5246_ack
      -- 
    phi_stmt_5246_ack_14438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_5246_ack_0, ack => zeropad3D_CP_2152_elements(1188)); -- 
    -- CP-element group 1189:  transition  input  bypass 
    -- CP-element group 1189: predecessors 
    -- CP-element group 1189: 	1187 
    -- CP-element group 1189: successors 
    -- CP-element group 1189: 	1191 
    -- CP-element group 1189:  members (1) 
      -- CP-element group 1189: 	 branch_block_stmt_714/merge_stmt_5245_PhiAck/phi_stmt_5253_ack
      -- 
    phi_stmt_5253_ack_14439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_5253_ack_0, ack => zeropad3D_CP_2152_elements(1189)); -- 
    -- CP-element group 1190:  transition  input  bypass 
    -- CP-element group 1190: predecessors 
    -- CP-element group 1190: 	1187 
    -- CP-element group 1190: successors 
    -- CP-element group 1190: 	1191 
    -- CP-element group 1190:  members (1) 
      -- CP-element group 1190: 	 branch_block_stmt_714/merge_stmt_5245_PhiAck/phi_stmt_5259_ack
      -- 
    phi_stmt_5259_ack_14440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_5259_ack_0, ack => zeropad3D_CP_2152_elements(1190)); -- 
    -- CP-element group 1191:  join  transition  bypass 
    -- CP-element group 1191: predecessors 
    -- CP-element group 1191: 	1188 
    -- CP-element group 1191: 	1189 
    -- CP-element group 1191: 	1190 
    -- CP-element group 1191: successors 
    -- CP-element group 1191: 	8 
    -- CP-element group 1191:  members (1) 
      -- CP-element group 1191: 	 branch_block_stmt_714/merge_stmt_5245_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_1191: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_cp_element_group_1191"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_2152_elements(1188) & zeropad3D_CP_2152_elements(1189) & zeropad3D_CP_2152_elements(1190);
      gj_zeropad3D_cp_element_group_1191 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_2152_elements(1191), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1059_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1143_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1168_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1393_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1408_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1432_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1458_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1616_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1699_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1724_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1945_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1960_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1984_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2010_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2174_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2257_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2282_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2520_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2535_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2559_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2585_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2742_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2825_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2850_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3071_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3086_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3110_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3136_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3306_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3389_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3414_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3658_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3673_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3697_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3723_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3886_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3969_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3994_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4227_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4242_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4266_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4292_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4450_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4533_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4558_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4796_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4811_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4835_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_4861_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_5012_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_5095_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_5120_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_829_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_844_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_868_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_894_wire : std_logic_vector(31 downto 0);
    signal LOAD_col_high_1234_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1234_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1331_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1331_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1555_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1555_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1790_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1790_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_1899_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_1899_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2107_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2107_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2348_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2348_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2445_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2445_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2681_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2681_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_2916_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_2916_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3025_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3025_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3239_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3239_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3480_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3480_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3583_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3583_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_3825_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_3825_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4060_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4060_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4181_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4181_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4383_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4383_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4624_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4624_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4715_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4715_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_4951_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_4951_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_5186_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_5186_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_782_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_782_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_col_high_992_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_col_high_992_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_1347_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_1347_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_1896_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_1896_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_2474_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_2474_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_3022_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_3022_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_3612_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_3612_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_4178_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_4178_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_4750_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_4750_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_depth_high_779_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_depth_high_779_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1344_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1344_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1893_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1893_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_2471_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2471_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3019_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3019_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3609_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3609_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_4175_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_4175_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_4747_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_4747_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_776_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_776_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1278_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1278_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1504_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1504_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1827_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1827_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_1880_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_1880_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2056_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2056_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2392_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2392_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2458_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2458_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2630_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2630_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_2953_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_2953_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3006_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3006_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3182_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3182_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3524_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3524_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3596_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3596_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_3768_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_3768_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4097_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4097_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4156_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4156_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4338_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4338_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4668_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4668_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4728_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4728_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_4906_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_4906_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_5223_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_5223_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_row_high_941_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_row_high_941_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom1002_3425_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1002_3425_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1177_3897_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1177_3897_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1220_3980_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1220_3980_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1225_4005_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1225_4005_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom130_1154_resized : std_logic_vector(13 downto 0);
    signal R_idxprom130_1154_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom135_1179_resized : std_logic_vector(13 downto 0);
    signal R_idxprom135_1179_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1395_4461_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1395_4461_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1438_4544_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1438_4544_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1443_4569_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1443_4569_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1615_5023_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1615_5023_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1658_5106_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1658_5106_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1663_5131_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1663_5131_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom298_1627_resized : std_logic_vector(13 downto 0);
    signal R_idxprom298_1627_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom341_1710_resized : std_logic_vector(13 downto 0);
    signal R_idxprom341_1710_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom346_1735_resized : std_logic_vector(13 downto 0);
    signal R_idxprom346_1735_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom515_2185_resized : std_logic_vector(13 downto 0);
    signal R_idxprom515_2185_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom558_2268_resized : std_logic_vector(13 downto 0);
    signal R_idxprom558_2268_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom563_2293_resized : std_logic_vector(13 downto 0);
    signal R_idxprom563_2293_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom736_2753_resized : std_logic_vector(13 downto 0);
    signal R_idxprom736_2753_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom779_2836_resized : std_logic_vector(13 downto 0);
    signal R_idxprom779_2836_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom784_2861_resized : std_logic_vector(13 downto 0);
    signal R_idxprom784_2861_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom954_3317_resized : std_logic_vector(13 downto 0);
    signal R_idxprom954_3317_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom997_3400_resized : std_logic_vector(13 downto 0);
    signal R_idxprom997_3400_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1071_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1071_scaled : std_logic_vector(13 downto 0);
    signal STORE_col_high_752_data_0 : std_logic_vector(7 downto 0);
    signal STORE_col_high_752_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_depth_high_771_data_0 : std_logic_vector(7 downto 0);
    signal STORE_depth_high_771_word_address_0 : std_logic_vector(0 downto 0);
    signal STORE_row_high_733_data_0 : std_logic_vector(7 downto 0);
    signal STORE_row_high_733_word_address_0 : std_logic_vector(0 downto 0);
    signal add1009_3445 : std_logic_vector(31 downto 0);
    signal add1017_3465 : std_logic_vector(15 downto 0);
    signal add102_1111 : std_logic_vector(31 downto 0);
    signal add1030_3496 : std_logic_vector(31 downto 0);
    signal add1047_3546 : std_logic_vector(31 downto 0);
    signal add111_1116 : std_logic_vector(31 downto 0);
    signal add1138_3790 : std_logic_vector(31 downto 0);
    signal add1155_3835 : std_logic_vector(31 downto 0);
    signal add1168_3874 : std_logic_vector(31 downto 0);
    signal add1174_3879 : std_logic_vector(31 downto 0);
    signal add1192_3937 : std_logic_vector(31 downto 0);
    signal add1201_3942 : std_logic_vector(31 downto 0);
    signal add1211_3957 : std_logic_vector(31 downto 0);
    signal add1217_3962 : std_logic_vector(31 downto 0);
    signal add121_1131 : std_logic_vector(31 downto 0);
    signal add1232_4025 : std_logic_vector(31 downto 0);
    signal add1240_4045 : std_logic_vector(15 downto 0);
    signal add1252_4070 : std_logic_vector(31 downto 0);
    signal add1269_4119 : std_logic_vector(31 downto 0);
    signal add127_1136 : std_logic_vector(31 downto 0);
    signal add1355_4348 : std_logic_vector(31 downto 0);
    signal add1373_4399 : std_logic_vector(31 downto 0);
    signal add1386_4438 : std_logic_vector(31 downto 0);
    signal add1392_4443 : std_logic_vector(31 downto 0);
    signal add140_1199 : std_logic_vector(31 downto 0);
    signal add1410_4501 : std_logic_vector(31 downto 0);
    signal add1419_4506 : std_logic_vector(31 downto 0);
    signal add1429_4521 : std_logic_vector(31 downto 0);
    signal add1435_4526 : std_logic_vector(31 downto 0);
    signal add1450_4589 : std_logic_vector(31 downto 0);
    signal add1458_4609 : std_logic_vector(15 downto 0);
    signal add1471_4640 : std_logic_vector(31 downto 0);
    signal add1486_4678 : std_logic_vector(31 downto 0);
    signal add148_1219 : std_logic_vector(15 downto 0);
    signal add1576_4916 : std_logic_vector(31 downto 0);
    signal add1593_4961 : std_logic_vector(31 downto 0);
    signal add159_1250 : std_logic_vector(31 downto 0);
    signal add1606_5000 : std_logic_vector(31 downto 0);
    signal add1612_5005 : std_logic_vector(31 downto 0);
    signal add1630_5063 : std_logic_vector(31 downto 0);
    signal add1639_5068 : std_logic_vector(31 downto 0);
    signal add1649_5083 : std_logic_vector(31 downto 0);
    signal add1655_5088 : std_logic_vector(31 downto 0);
    signal add1670_5151 : std_logic_vector(31 downto 0);
    signal add1678_5171 : std_logic_vector(15 downto 0);
    signal add1690_5196 : std_logic_vector(31 downto 0);
    signal add1705_5233 : std_logic_vector(31 downto 0);
    signal add175_1294 : std_logic_vector(31 downto 0);
    signal add259_1520 : std_logic_vector(31 downto 0);
    signal add276_1565 : std_logic_vector(31 downto 0);
    signal add289_1604 : std_logic_vector(31 downto 0);
    signal add295_1609 : std_logic_vector(31 downto 0);
    signal add313_1667 : std_logic_vector(31 downto 0);
    signal add322_1672 : std_logic_vector(31 downto 0);
    signal add332_1687 : std_logic_vector(31 downto 0);
    signal add338_1692 : std_logic_vector(31 downto 0);
    signal add353_1755 : std_logic_vector(31 downto 0);
    signal add361_1775 : std_logic_vector(15 downto 0);
    signal add373_1800 : std_logic_vector(31 downto 0);
    signal add389_1843 : std_logic_vector(31 downto 0);
    signal add475_2072 : std_logic_vector(31 downto 0);
    signal add493_2123 : std_logic_vector(31 downto 0);
    signal add506_2162 : std_logic_vector(31 downto 0);
    signal add512_2167 : std_logic_vector(31 downto 0);
    signal add530_2225 : std_logic_vector(31 downto 0);
    signal add539_2230 : std_logic_vector(31 downto 0);
    signal add549_2245 : std_logic_vector(31 downto 0);
    signal add555_2250 : std_logic_vector(31 downto 0);
    signal add570_2313 : std_logic_vector(31 downto 0);
    signal add578_2333 : std_logic_vector(15 downto 0);
    signal add591_2364 : std_logic_vector(31 downto 0);
    signal add607_2408 : std_logic_vector(31 downto 0);
    signal add697_2646 : std_logic_vector(31 downto 0);
    signal add714_2691 : std_logic_vector(31 downto 0);
    signal add727_2730 : std_logic_vector(31 downto 0);
    signal add733_2735 : std_logic_vector(31 downto 0);
    signal add73_1008 : std_logic_vector(31 downto 0);
    signal add751_2793 : std_logic_vector(31 downto 0);
    signal add760_2798 : std_logic_vector(31 downto 0);
    signal add770_2813 : std_logic_vector(31 downto 0);
    signal add776_2818 : std_logic_vector(31 downto 0);
    signal add791_2881 : std_logic_vector(31 downto 0);
    signal add799_2901 : std_logic_vector(15 downto 0);
    signal add811_2926 : std_logic_vector(31 downto 0);
    signal add827_2969 : std_logic_vector(31 downto 0);
    signal add84_1047 : std_logic_vector(31 downto 0);
    signal add90_1052 : std_logic_vector(31 downto 0);
    signal add914_3204 : std_logic_vector(31 downto 0);
    signal add932_3255 : std_logic_vector(31 downto 0);
    signal add945_3294 : std_logic_vector(31 downto 0);
    signal add951_3299 : std_logic_vector(31 downto 0);
    signal add969_3357 : std_logic_vector(31 downto 0);
    signal add978_3362 : std_logic_vector(31 downto 0);
    signal add988_3377 : std_logic_vector(31 downto 0);
    signal add994_3382 : std_logic_vector(31 downto 0);
    signal add_957 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1072_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1155_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1180_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1628_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1628_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1628_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1628_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1628_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1628_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1711_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1736_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2186_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2186_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2186_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2186_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2186_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2186_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2269_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2269_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2269_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2269_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2269_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2269_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2294_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2294_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2294_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2294_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2294_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2294_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2754_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2754_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2754_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2754_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2754_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2754_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2837_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2837_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2837_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2837_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2837_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2837_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2862_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2862_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2862_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2862_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2862_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2862_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3318_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3318_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3318_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3318_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3318_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3318_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3401_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3401_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3401_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3401_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3401_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3401_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3426_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3426_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3426_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3426_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3426_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3426_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3898_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3898_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3898_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3898_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3898_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3898_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3981_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3981_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3981_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3981_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3981_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3981_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4006_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4006_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4006_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4006_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4006_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4006_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4462_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4462_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4462_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4462_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4462_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4462_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4545_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4545_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4545_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4545_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4545_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4545_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4570_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4570_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_4570_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4570_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_4570_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_4570_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5024_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5024_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5024_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5024_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5024_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5024_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5107_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5107_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5107_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5107_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5107_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5107_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5132_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5132_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_5132_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5132_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_5132_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_5132_root_address : std_logic_vector(13 downto 0);
    signal arrayidx1003_3428 : std_logic_vector(31 downto 0);
    signal arrayidx1178_3900 : std_logic_vector(31 downto 0);
    signal arrayidx1221_3983 : std_logic_vector(31 downto 0);
    signal arrayidx1226_4008 : std_logic_vector(31 downto 0);
    signal arrayidx131_1157 : std_logic_vector(31 downto 0);
    signal arrayidx136_1182 : std_logic_vector(31 downto 0);
    signal arrayidx1396_4464 : std_logic_vector(31 downto 0);
    signal arrayidx1439_4547 : std_logic_vector(31 downto 0);
    signal arrayidx1444_4572 : std_logic_vector(31 downto 0);
    signal arrayidx1616_5026 : std_logic_vector(31 downto 0);
    signal arrayidx1659_5109 : std_logic_vector(31 downto 0);
    signal arrayidx1664_5134 : std_logic_vector(31 downto 0);
    signal arrayidx299_1630 : std_logic_vector(31 downto 0);
    signal arrayidx342_1713 : std_logic_vector(31 downto 0);
    signal arrayidx347_1738 : std_logic_vector(31 downto 0);
    signal arrayidx516_2188 : std_logic_vector(31 downto 0);
    signal arrayidx559_2271 : std_logic_vector(31 downto 0);
    signal arrayidx564_2296 : std_logic_vector(31 downto 0);
    signal arrayidx737_2756 : std_logic_vector(31 downto 0);
    signal arrayidx780_2839 : std_logic_vector(31 downto 0);
    signal arrayidx785_2864 : std_logic_vector(31 downto 0);
    signal arrayidx955_3320 : std_logic_vector(31 downto 0);
    signal arrayidx998_3403 : std_logic_vector(31 downto 0);
    signal arrayidx_1074 : std_logic_vector(31 downto 0);
    signal call_716 : std_logic_vector(15 downto 0);
    signal cmp1012_3452 : std_logic_vector(0 downto 0);
    signal cmp1031_3501 : std_logic_vector(0 downto 0);
    signal cmp1048_3551 : std_logic_vector(0 downto 0);
    signal cmp1127_3759 : std_logic_vector(0 downto 0);
    signal cmp1139_3797 : std_logic_vector(0 downto 0);
    signal cmp1146_3816 : std_logic_vector(0 downto 0);
    signal cmp1156_3842 : std_logic_vector(0 downto 0);
    signal cmp1235_4032 : std_logic_vector(0 downto 0);
    signal cmp1253_4075 : std_logic_vector(0 downto 0);
    signal cmp1270_4124 : std_logic_vector(0 downto 0);
    signal cmp1346_4329 : std_logic_vector(0 downto 0);
    signal cmp1356_4355 : std_logic_vector(0 downto 0);
    signal cmp1363_4374 : std_logic_vector(0 downto 0);
    signal cmp1374_4406 : std_logic_vector(0 downto 0);
    signal cmp143_1206 : std_logic_vector(0 downto 0);
    signal cmp1453_4596 : std_logic_vector(0 downto 0);
    signal cmp1472_4645 : std_logic_vector(0 downto 0);
    signal cmp1487_4683 : std_logic_vector(0 downto 0);
    signal cmp1567_4897 : std_logic_vector(0 downto 0);
    signal cmp1577_4923 : std_logic_vector(0 downto 0);
    signal cmp1584_4942 : std_logic_vector(0 downto 0);
    signal cmp1594_4968 : std_logic_vector(0 downto 0);
    signal cmp160_1255 : std_logic_vector(0 downto 0);
    signal cmp1673_5158 : std_logic_vector(0 downto 0);
    signal cmp1691_5201 : std_logic_vector(0 downto 0);
    signal cmp1706_5238 : std_logic_vector(0 downto 0);
    signal cmp176_1299 : std_logic_vector(0 downto 0);
    signal cmp249_1495 : std_logic_vector(0 downto 0);
    signal cmp260_1527 : std_logic_vector(0 downto 0);
    signal cmp267_1546 : std_logic_vector(0 downto 0);
    signal cmp277_1572 : std_logic_vector(0 downto 0);
    signal cmp356_1762 : std_logic_vector(0 downto 0);
    signal cmp374_1805 : std_logic_vector(0 downto 0);
    signal cmp390_1848 : std_logic_vector(0 downto 0);
    signal cmp465_2047 : std_logic_vector(0 downto 0);
    signal cmp476_2079 : std_logic_vector(0 downto 0);
    signal cmp483_2098 : std_logic_vector(0 downto 0);
    signal cmp494_2130 : std_logic_vector(0 downto 0);
    signal cmp56_964 : std_logic_vector(0 downto 0);
    signal cmp573_2320 : std_logic_vector(0 downto 0);
    signal cmp592_2369 : std_logic_vector(0 downto 0);
    signal cmp608_2413 : std_logic_vector(0 downto 0);
    signal cmp63_983 : std_logic_vector(0 downto 0);
    signal cmp687_2621 : std_logic_vector(0 downto 0);
    signal cmp698_2653 : std_logic_vector(0 downto 0);
    signal cmp705_2672 : std_logic_vector(0 downto 0);
    signal cmp715_2698 : std_logic_vector(0 downto 0);
    signal cmp74_1015 : std_logic_vector(0 downto 0);
    signal cmp794_2888 : std_logic_vector(0 downto 0);
    signal cmp812_2931 : std_logic_vector(0 downto 0);
    signal cmp828_2974 : std_logic_vector(0 downto 0);
    signal cmp903_3173 : std_logic_vector(0 downto 0);
    signal cmp915_3211 : std_logic_vector(0 downto 0);
    signal cmp922_3230 : std_logic_vector(0 downto 0);
    signal cmp933_3262 : std_logic_vector(0 downto 0);
    signal cmp_932 : std_logic_vector(0 downto 0);
    signal conv1008_3439 : std_logic_vector(31 downto 0);
    signal conv1023_3478 : std_logic_vector(31 downto 0);
    signal conv1025_3485 : std_logic_vector(31 downto 0);
    signal conv1039_3522 : std_logic_vector(31 downto 0);
    signal conv1041_3529 : std_logic_vector(31 downto 0);
    signal conv104_896 : std_logic_vector(31 downto 0);
    signal conv1064_3588 : std_logic_vector(15 downto 0);
    signal conv1070_3601 : std_logic_vector(15 downto 0);
    signal conv1104_3641 : std_logic_vector(31 downto 0);
    signal conv1106_3645 : std_logic_vector(31 downto 0);
    signal conv1112_3660 : std_logic_vector(31 downto 0);
    signal conv1114_3675 : std_logic_vector(31 downto 0);
    signal conv1124_3752 : std_logic_vector(31 downto 0);
    signal conv1126_3684 : std_logic_vector(31 downto 0);
    signal conv1133_3773 : std_logic_vector(31 downto 0);
    signal conv1143_3809 : std_logic_vector(31 downto 0);
    signal conv1152_3830 : std_logic_vector(31 downto 0);
    signal conv1162_3854 : std_logic_vector(31 downto 0);
    signal conv1166_3859 : std_logic_vector(31 downto 0);
    signal conv1170_3699 : std_logic_vector(31 downto 0);
    signal conv1183_3912 : std_logic_vector(31 downto 0);
    signal conv1194_3725 : std_logic_vector(31 downto 0);
    signal conv1231_4019 : std_logic_vector(31 downto 0);
    signal conv1246_4058 : std_logic_vector(31 downto 0);
    signal conv1248_4065 : std_logic_vector(31 downto 0);
    signal conv1261_4095 : std_logic_vector(31 downto 0);
    signal conv1263_4102 : std_logic_vector(31 downto 0);
    signal conv1288_4161 : std_logic_vector(15 downto 0);
    signal conv1323_4210 : std_logic_vector(31 downto 0);
    signal conv1325_4214 : std_logic_vector(31 downto 0);
    signal conv1331_4229 : std_logic_vector(31 downto 0);
    signal conv1333_4244 : std_logic_vector(31 downto 0);
    signal conv1343_4322 : std_logic_vector(31 downto 0);
    signal conv1345_4253 : std_logic_vector(31 downto 0);
    signal conv1352_4343 : std_logic_vector(31 downto 0);
    signal conv1360_4367 : std_logic_vector(31 downto 0);
    signal conv1369_4388 : std_logic_vector(31 downto 0);
    signal conv1380_4418 : std_logic_vector(31 downto 0);
    signal conv1384_4423 : std_logic_vector(31 downto 0);
    signal conv1388_4268 : std_logic_vector(31 downto 0);
    signal conv139_1193 : std_logic_vector(31 downto 0);
    signal conv1401_4476 : std_logic_vector(31 downto 0);
    signal conv1412_4294 : std_logic_vector(31 downto 0);
    signal conv1449_4583 : std_logic_vector(31 downto 0);
    signal conv1464_4622 : std_logic_vector(31 downto 0);
    signal conv1466_4629 : std_logic_vector(31 downto 0);
    signal conv1480_4666 : std_logic_vector(31 downto 0);
    signal conv1482_4673 : std_logic_vector(31 downto 0);
    signal conv1503_4720 : std_logic_vector(15 downto 0);
    signal conv1509_4733 : std_logic_vector(15 downto 0);
    signal conv153_1232 : std_logic_vector(31 downto 0);
    signal conv1544_4779 : std_logic_vector(31 downto 0);
    signal conv1546_4783 : std_logic_vector(31 downto 0);
    signal conv1552_4798 : std_logic_vector(31 downto 0);
    signal conv1554_4813 : std_logic_vector(31 downto 0);
    signal conv155_1239 : std_logic_vector(31 downto 0);
    signal conv1564_4890 : std_logic_vector(31 downto 0);
    signal conv1566_4822 : std_logic_vector(31 downto 0);
    signal conv1573_4911 : std_logic_vector(31 downto 0);
    signal conv1581_4935 : std_logic_vector(31 downto 0);
    signal conv1590_4956 : std_logic_vector(31 downto 0);
    signal conv1600_4980 : std_logic_vector(31 downto 0);
    signal conv1604_4985 : std_logic_vector(31 downto 0);
    signal conv1608_4837 : std_logic_vector(31 downto 0);
    signal conv1621_5038 : std_logic_vector(31 downto 0);
    signal conv1632_4863 : std_logic_vector(31 downto 0);
    signal conv1669_5145 : std_logic_vector(31 downto 0);
    signal conv1684_5184 : std_logic_vector(31 downto 0);
    signal conv1686_5191 : std_logic_vector(31 downto 0);
    signal conv168_1276 : std_logic_vector(31 downto 0);
    signal conv1699_5221 : std_logic_vector(31 downto 0);
    signal conv1701_5228 : std_logic_vector(31 downto 0);
    signal conv170_1283 : std_logic_vector(31 downto 0);
    signal conv190_1336 : std_logic_vector(15 downto 0);
    signal conv226_1376 : std_logic_vector(31 downto 0);
    signal conv228_1380 : std_logic_vector(31 downto 0);
    signal conv234_1395 : std_logic_vector(31 downto 0);
    signal conv236_1410 : std_logic_vector(31 downto 0);
    signal conv246_1488 : std_logic_vector(31 downto 0);
    signal conv248_1419 : std_logic_vector(31 downto 0);
    signal conv255_1509 : std_logic_vector(31 downto 0);
    signal conv264_1539 : std_logic_vector(31 downto 0);
    signal conv273_1560 : std_logic_vector(31 downto 0);
    signal conv283_1584 : std_logic_vector(31 downto 0);
    signal conv287_1589 : std_logic_vector(31 downto 0);
    signal conv291_1434 : std_logic_vector(31 downto 0);
    signal conv2_751 : std_logic_vector(7 downto 0);
    signal conv304_1642 : std_logic_vector(31 downto 0);
    signal conv315_1460 : std_logic_vector(31 downto 0);
    signal conv31_811 : std_logic_vector(31 downto 0);
    signal conv33_815 : std_logic_vector(31 downto 0);
    signal conv352_1749 : std_logic_vector(31 downto 0);
    signal conv367_1788 : std_logic_vector(31 downto 0);
    signal conv369_1795 : std_logic_vector(31 downto 0);
    signal conv37_831 : std_logic_vector(31 downto 0);
    signal conv382_1825 : std_logic_vector(31 downto 0);
    signal conv384_1832 : std_logic_vector(31 downto 0);
    signal conv39_846 : std_logic_vector(31 downto 0);
    signal conv408_1885 : std_logic_vector(15 downto 0);
    signal conv442_1928 : std_logic_vector(31 downto 0);
    signal conv444_1932 : std_logic_vector(31 downto 0);
    signal conv450_1947 : std_logic_vector(31 downto 0);
    signal conv452_1962 : std_logic_vector(31 downto 0);
    signal conv462_2040 : std_logic_vector(31 downto 0);
    signal conv464_1971 : std_logic_vector(31 downto 0);
    signal conv46_925 : std_logic_vector(31 downto 0);
    signal conv471_2061 : std_logic_vector(31 downto 0);
    signal conv480_2091 : std_logic_vector(31 downto 0);
    signal conv489_2112 : std_logic_vector(31 downto 0);
    signal conv48_855 : std_logic_vector(31 downto 0);
    signal conv4_770 : std_logic_vector(7 downto 0);
    signal conv500_2142 : std_logic_vector(31 downto 0);
    signal conv504_2147 : std_logic_vector(31 downto 0);
    signal conv508_1986 : std_logic_vector(31 downto 0);
    signal conv521_2200 : std_logic_vector(31 downto 0);
    signal conv532_2012 : std_logic_vector(31 downto 0);
    signal conv53_946 : std_logic_vector(31 downto 0);
    signal conv569_2307 : std_logic_vector(31 downto 0);
    signal conv584_2346 : std_logic_vector(31 downto 0);
    signal conv586_2353 : std_logic_vector(31 downto 0);
    signal conv600_2390 : std_logic_vector(31 downto 0);
    signal conv602_2397 : std_logic_vector(31 downto 0);
    signal conv60_976 : std_logic_vector(31 downto 0);
    signal conv624_2450 : std_logic_vector(15 downto 0);
    signal conv630_2463 : std_logic_vector(15 downto 0);
    signal conv664_2503 : std_logic_vector(31 downto 0);
    signal conv666_2507 : std_logic_vector(31 downto 0);
    signal conv672_2522 : std_logic_vector(31 downto 0);
    signal conv674_2537 : std_logic_vector(31 downto 0);
    signal conv684_2614 : std_logic_vector(31 downto 0);
    signal conv686_2546 : std_logic_vector(31 downto 0);
    signal conv693_2635 : std_logic_vector(31 downto 0);
    signal conv69_997 : std_logic_vector(31 downto 0);
    signal conv702_2665 : std_logic_vector(31 downto 0);
    signal conv711_2686 : std_logic_vector(31 downto 0);
    signal conv721_2710 : std_logic_vector(31 downto 0);
    signal conv725_2715 : std_logic_vector(31 downto 0);
    signal conv729_2561 : std_logic_vector(31 downto 0);
    signal conv742_2768 : std_logic_vector(31 downto 0);
    signal conv753_2587 : std_logic_vector(31 downto 0);
    signal conv78_1027 : std_logic_vector(31 downto 0);
    signal conv790_2875 : std_logic_vector(31 downto 0);
    signal conv805_2914 : std_logic_vector(31 downto 0);
    signal conv807_2921 : std_logic_vector(31 downto 0);
    signal conv820_2951 : std_logic_vector(31 downto 0);
    signal conv822_2958 : std_logic_vector(31 downto 0);
    signal conv82_1032 : std_logic_vector(31 downto 0);
    signal conv846_3011 : std_logic_vector(15 downto 0);
    signal conv86_870 : std_logic_vector(31 downto 0);
    signal conv880_3054 : std_logic_vector(31 downto 0);
    signal conv882_3058 : std_logic_vector(31 downto 0);
    signal conv888_3073 : std_logic_vector(31 downto 0);
    signal conv890_3088 : std_logic_vector(31 downto 0);
    signal conv900_3166 : std_logic_vector(31 downto 0);
    signal conv902_3097 : std_logic_vector(31 downto 0);
    signal conv909_3187 : std_logic_vector(31 downto 0);
    signal conv919_3223 : std_logic_vector(31 downto 0);
    signal conv928_3244 : std_logic_vector(31 downto 0);
    signal conv939_3274 : std_logic_vector(31 downto 0);
    signal conv943_3279 : std_logic_vector(31 downto 0);
    signal conv947_3112 : std_logic_vector(31 downto 0);
    signal conv94_1086 : std_logic_vector(31 downto 0);
    signal conv960_3332 : std_logic_vector(31 downto 0);
    signal conv971_3138 : std_logic_vector(31 downto 0);
    signal conv_732 : std_logic_vector(7 downto 0);
    signal div1026_3491 : std_logic_vector(31 downto 0);
    signal div1043_3541 : std_logic_vector(31 downto 0);
    signal div1065_3594 : std_logic_vector(15 downto 0);
    signal div1071_3607 : std_logic_vector(15 downto 0);
    signal div1135_3785 : std_logic_vector(31 downto 0);
    signal div1265_4114 : std_logic_vector(31 downto 0);
    signal div1289_4167 : std_logic_vector(15 downto 0);
    signal div1370_4394 : std_logic_vector(31 downto 0);
    signal div1467_4635 : std_logic_vector(31 downto 0);
    signal div1504_4726 : std_logic_vector(15 downto 0);
    signal div1511_4745 : std_logic_vector(15 downto 0);
    signal div156_1245 : std_logic_vector(31 downto 0);
    signal div171_1289 : std_logic_vector(31 downto 0);
    signal div191_1342 : std_logic_vector(15 downto 0);
    signal div256_1515 : std_logic_vector(31 downto 0);
    signal div385_1838 : std_logic_vector(31 downto 0);
    signal div409_1891 : std_logic_vector(15 downto 0);
    signal div472_2067 : std_logic_vector(31 downto 0);
    signal div490_2118 : std_logic_vector(31 downto 0);
    signal div587_2359 : std_logic_vector(31 downto 0);
    signal div603_2403 : std_logic_vector(31 downto 0);
    signal div625_2456 : std_logic_vector(15 downto 0);
    signal div631_2469 : std_logic_vector(15 downto 0);
    signal div694_2641 : std_logic_vector(31 downto 0);
    signal div70_1003 : std_logic_vector(31 downto 0);
    signal div823_2964 : std_logic_vector(31 downto 0);
    signal div847_3017 : std_logic_vector(15 downto 0);
    signal div911_3199 : std_logic_vector(31 downto 0);
    signal div929_3250 : std_logic_vector(31 downto 0);
    signal div_952 : std_logic_vector(31 downto 0);
    signal i1068x_x1x_xph_4139 : std_logic_vector(15 downto 0);
    signal i1068x_x2_3735 : std_logic_vector(15 downto 0);
    signal i1286x_x1x_xph_4698 : std_logic_vector(15 downto 0);
    signal i1286x_x2_4304 : std_logic_vector(15 downto 0);
    signal i1507x_x1x_xph_5253 : std_logic_vector(15 downto 0);
    signal i1507x_x2_4873 : std_logic_vector(15 downto 0);
    signal i194x_x1x_xph_1862 : std_logic_vector(15 downto 0);
    signal i194x_x2_1469 : std_logic_vector(15 downto 0);
    signal i406x_x1x_xph_2428 : std_logic_vector(15 downto 0);
    signal i406x_x2_2022 : std_logic_vector(15 downto 0);
    signal i628x_x1x_xph_2989 : std_logic_vector(15 downto 0);
    signal i628x_x2_2597 : std_logic_vector(15 downto 0);
    signal i844x_x1x_xph_3566 : std_logic_vector(15 downto 0);
    signal i844x_x2_3148 : std_logic_vector(15 downto 0);
    signal iNsTr_0_724 : std_logic_vector(31 downto 0);
    signal iNsTr_107_4190 : std_logic_vector(31 downto 0);
    signal iNsTr_108_4202 : std_logic_vector(31 downto 0);
    signal iNsTr_124_4759 : std_logic_vector(31 downto 0);
    signal iNsTr_125_4771 : std_logic_vector(31 downto 0);
    signal iNsTr_22_1356 : std_logic_vector(31 downto 0);
    signal iNsTr_23_1368 : std_logic_vector(31 downto 0);
    signal iNsTr_2_743 : std_logic_vector(31 downto 0);
    signal iNsTr_39_1908 : std_logic_vector(31 downto 0);
    signal iNsTr_40_1920 : std_logic_vector(31 downto 0);
    signal iNsTr_4_762 : std_logic_vector(31 downto 0);
    signal iNsTr_56_2483 : std_logic_vector(31 downto 0);
    signal iNsTr_57_2495 : std_logic_vector(31 downto 0);
    signal iNsTr_73_3034 : std_logic_vector(31 downto 0);
    signal iNsTr_74_3046 : std_logic_vector(31 downto 0);
    signal iNsTr_7_791 : std_logic_vector(31 downto 0);
    signal iNsTr_8_803 : std_logic_vector(31 downto 0);
    signal iNsTr_90_3621 : std_logic_vector(31 downto 0);
    signal iNsTr_91_3633 : std_logic_vector(31 downto 0);
    signal idxprom1002_3421 : std_logic_vector(63 downto 0);
    signal idxprom1177_3893 : std_logic_vector(63 downto 0);
    signal idxprom1220_3976 : std_logic_vector(63 downto 0);
    signal idxprom1225_4001 : std_logic_vector(63 downto 0);
    signal idxprom130_1150 : std_logic_vector(63 downto 0);
    signal idxprom135_1175 : std_logic_vector(63 downto 0);
    signal idxprom1395_4457 : std_logic_vector(63 downto 0);
    signal idxprom1438_4540 : std_logic_vector(63 downto 0);
    signal idxprom1443_4565 : std_logic_vector(63 downto 0);
    signal idxprom1615_5019 : std_logic_vector(63 downto 0);
    signal idxprom1658_5102 : std_logic_vector(63 downto 0);
    signal idxprom1663_5127 : std_logic_vector(63 downto 0);
    signal idxprom298_1623 : std_logic_vector(63 downto 0);
    signal idxprom341_1706 : std_logic_vector(63 downto 0);
    signal idxprom346_1731 : std_logic_vector(63 downto 0);
    signal idxprom515_2181 : std_logic_vector(63 downto 0);
    signal idxprom558_2264 : std_logic_vector(63 downto 0);
    signal idxprom563_2289 : std_logic_vector(63 downto 0);
    signal idxprom736_2749 : std_logic_vector(63 downto 0);
    signal idxprom779_2832 : std_logic_vector(63 downto 0);
    signal idxprom784_2857 : std_logic_vector(63 downto 0);
    signal idxprom954_3313 : std_logic_vector(63 downto 0);
    signal idxprom997_3396 : std_logic_vector(63 downto 0);
    signal idxprom_1067 : std_logic_vector(63 downto 0);
    signal inc1021_3473 : std_logic_vector(15 downto 0);
    signal inc1036_3505 : std_logic_vector(15 downto 0);
    signal inc1036x_xi844x_x2_3510 : std_logic_vector(15 downto 0);
    signal inc1244_4053 : std_logic_vector(15 downto 0);
    signal inc1258_4079 : std_logic_vector(15 downto 0);
    signal inc1258x_xi1068x_x2_4084 : std_logic_vector(15 downto 0);
    signal inc1462_4617 : std_logic_vector(15 downto 0);
    signal inc1477_4649 : std_logic_vector(15 downto 0);
    signal inc1477x_xi1286x_x2_4654 : std_logic_vector(15 downto 0);
    signal inc165_1259 : std_logic_vector(15 downto 0);
    signal inc165x_xix_x2_1264 : std_logic_vector(15 downto 0);
    signal inc1682_5179 : std_logic_vector(15 downto 0);
    signal inc1696_5205 : std_logic_vector(15 downto 0);
    signal inc1696x_xi1507x_x2_5210 : std_logic_vector(15 downto 0);
    signal inc365_1783 : std_logic_vector(15 downto 0);
    signal inc379_1809 : std_logic_vector(15 downto 0);
    signal inc379x_xi194x_x2_1814 : std_logic_vector(15 downto 0);
    signal inc582_2341 : std_logic_vector(15 downto 0);
    signal inc597_2373 : std_logic_vector(15 downto 0);
    signal inc597x_xi406x_x2_2378 : std_logic_vector(15 downto 0);
    signal inc803_2909 : std_logic_vector(15 downto 0);
    signal inc817_2935 : std_logic_vector(15 downto 0);
    signal inc817x_xi628x_x2_2940 : std_logic_vector(15 downto 0);
    signal inc_1227 : std_logic_vector(15 downto 0);
    signal ix_x1x_xph_1313 : std_logic_vector(15 downto 0);
    signal ix_x2_906 : std_logic_vector(15 downto 0);
    signal j1118x_x0x_xph_4145 : std_logic_vector(15 downto 0);
    signal j1118x_x1_3741 : std_logic_vector(15 downto 0);
    signal j1118x_x2_4090 : std_logic_vector(15 downto 0);
    signal j1337x_x0x_xph_4704 : std_logic_vector(15 downto 0);
    signal j1337x_x1_4310 : std_logic_vector(15 downto 0);
    signal j1337x_x2_4661 : std_logic_vector(15 downto 0);
    signal j1558x_x0x_xph_5259 : std_logic_vector(15 downto 0);
    signal j1558x_x1_4879 : std_logic_vector(15 downto 0);
    signal j1558x_x2_5216 : std_logic_vector(15 downto 0);
    signal j240x_x0x_xph_1856 : std_logic_vector(15 downto 0);
    signal j240x_x1_1463 : std_logic_vector(15 downto 0);
    signal j240x_x2_1820 : std_logic_vector(15 downto 0);
    signal j456x_x0x_xph_2434 : std_logic_vector(15 downto 0);
    signal j456x_x1_2028 : std_logic_vector(15 downto 0);
    signal j456x_x2_2385 : std_logic_vector(15 downto 0);
    signal j678x_x0x_xph_2995 : std_logic_vector(15 downto 0);
    signal j678x_x1_2603 : std_logic_vector(15 downto 0);
    signal j678x_x2_2946 : std_logic_vector(15 downto 0);
    signal j894x_x0x_xph_3572 : std_logic_vector(15 downto 0);
    signal j894x_x1_3154 : std_logic_vector(15 downto 0);
    signal j894x_x2_3517 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_1307 : std_logic_vector(15 downto 0);
    signal jx_x1_899 : std_logic_vector(15 downto 0);
    signal jx_x2_1271 : std_logic_vector(15 downto 0);
    signal k1060x_x0x_xph_4132 : std_logic_vector(15 downto 0);
    signal k1060x_x1_3728 : std_logic_vector(15 downto 0);
    signal k1282x_x0x_xph_4691 : std_logic_vector(15 downto 0);
    signal k1282x_x1_4297 : std_logic_vector(15 downto 0);
    signal k1499x_x0x_xph_5246 : std_logic_vector(15 downto 0);
    signal k1499x_x1_4866 : std_logic_vector(15 downto 0);
    signal k186x_x0x_xph_1868 : std_logic_vector(15 downto 0);
    signal k186x_x1_1476 : std_logic_vector(15 downto 0);
    signal k402x_x0x_xph_2421 : std_logic_vector(15 downto 0);
    signal k402x_x1_2015 : std_logic_vector(15 downto 0);
    signal k620x_x0x_xph_2982 : std_logic_vector(15 downto 0);
    signal k620x_x1_2590 : std_logic_vector(15 downto 0);
    signal k840x_x0x_xph_3559 : std_logic_vector(15 downto 0);
    signal k840x_x1_3141 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_1319 : std_logic_vector(15 downto 0);
    signal kx_x1_913 : std_logic_vector(15 downto 0);
    signal mul101_1096 : std_logic_vector(31 downto 0);
    signal mul1042_3535 : std_logic_vector(31 downto 0);
    signal mul1107_3711 : std_logic_vector(31 downto 0);
    signal mul110_1106 : std_logic_vector(31 downto 0);
    signal mul1115_3680 : std_logic_vector(31 downto 0);
    signal mul1134_3779 : std_logic_vector(31 downto 0);
    signal mul1167_3864 : std_logic_vector(31 downto 0);
    signal mul1173_3869 : std_logic_vector(31 downto 0);
    signal mul1191_3922 : std_logic_vector(31 downto 0);
    signal mul1200_3932 : std_logic_vector(31 downto 0);
    signal mul120_1121 : std_logic_vector(31 downto 0);
    signal mul1210_3947 : std_logic_vector(31 downto 0);
    signal mul1216_3952 : std_logic_vector(31 downto 0);
    signal mul1264_4108 : std_logic_vector(31 downto 0);
    signal mul126_1126 : std_logic_vector(31 downto 0);
    signal mul1290_4173 : std_logic_vector(15 downto 0);
    signal mul1326_4280 : std_logic_vector(31 downto 0);
    signal mul1334_4249 : std_logic_vector(31 downto 0);
    signal mul1385_4428 : std_logic_vector(31 downto 0);
    signal mul1391_4433 : std_logic_vector(31 downto 0);
    signal mul1409_4486 : std_logic_vector(31 downto 0);
    signal mul1418_4496 : std_logic_vector(31 downto 0);
    signal mul1428_4511 : std_logic_vector(31 downto 0);
    signal mul1434_4516 : std_logic_vector(31 downto 0);
    signal mul1510_4739 : std_logic_vector(15 downto 0);
    signal mul1547_4849 : std_logic_vector(31 downto 0);
    signal mul1555_4818 : std_logic_vector(31 downto 0);
    signal mul1605_4990 : std_logic_vector(31 downto 0);
    signal mul1611_4995 : std_logic_vector(31 downto 0);
    signal mul1629_5048 : std_logic_vector(31 downto 0);
    signal mul1638_5058 : std_logic_vector(31 downto 0);
    signal mul1648_5073 : std_logic_vector(31 downto 0);
    signal mul1654_5078 : std_logic_vector(31 downto 0);
    signal mul229_1446 : std_logic_vector(31 downto 0);
    signal mul237_1415 : std_logic_vector(31 downto 0);
    signal mul288_1594 : std_logic_vector(31 downto 0);
    signal mul294_1599 : std_logic_vector(31 downto 0);
    signal mul312_1652 : std_logic_vector(31 downto 0);
    signal mul321_1662 : std_logic_vector(31 downto 0);
    signal mul331_1677 : std_logic_vector(31 downto 0);
    signal mul337_1682 : std_logic_vector(31 downto 0);
    signal mul40_851 : std_logic_vector(31 downto 0);
    signal mul445_1998 : std_logic_vector(31 downto 0);
    signal mul453_1967 : std_logic_vector(31 downto 0);
    signal mul505_2152 : std_logic_vector(31 downto 0);
    signal mul511_2157 : std_logic_vector(31 downto 0);
    signal mul529_2210 : std_logic_vector(31 downto 0);
    signal mul538_2220 : std_logic_vector(31 downto 0);
    signal mul548_2235 : std_logic_vector(31 downto 0);
    signal mul554_2240 : std_logic_vector(31 downto 0);
    signal mul667_2573 : std_logic_vector(31 downto 0);
    signal mul675_2542 : std_logic_vector(31 downto 0);
    signal mul726_2720 : std_logic_vector(31 downto 0);
    signal mul732_2725 : std_logic_vector(31 downto 0);
    signal mul750_2778 : std_logic_vector(31 downto 0);
    signal mul759_2788 : std_logic_vector(31 downto 0);
    signal mul769_2803 : std_logic_vector(31 downto 0);
    signal mul775_2808 : std_logic_vector(31 downto 0);
    signal mul83_1037 : std_logic_vector(31 downto 0);
    signal mul883_3124 : std_logic_vector(31 downto 0);
    signal mul891_3093 : std_logic_vector(31 downto 0);
    signal mul89_1042 : std_logic_vector(31 downto 0);
    signal mul910_3193 : std_logic_vector(31 downto 0);
    signal mul944_3284 : std_logic_vector(31 downto 0);
    signal mul950_3289 : std_logic_vector(31 downto 0);
    signal mul968_3342 : std_logic_vector(31 downto 0);
    signal mul977_3352 : std_logic_vector(31 downto 0);
    signal mul987_3367 : std_logic_vector(31 downto 0);
    signal mul993_3372 : std_logic_vector(31 downto 0);
    signal mul_882 : std_logic_vector(31 downto 0);
    signal ptr_deref_1076_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1076_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1076_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1076_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1160_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1160_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1184_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1184_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1184_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1359_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1359_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1371_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1371_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1371_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1371_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1371_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1632_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1632_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1632_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1632_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1632_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1632_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1716_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1716_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1740_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1740_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1740_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1911_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1911_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1911_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1911_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1911_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1923_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1923_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1923_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1923_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1923_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2190_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2190_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2190_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2190_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2190_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2190_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2274_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2274_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2274_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2274_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2274_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2298_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2298_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2298_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2298_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2298_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2298_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2486_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2486_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2486_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2486_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2486_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2498_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2758_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2758_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2758_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2758_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2758_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2758_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2842_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2842_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2842_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2842_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2842_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2866_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2866_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2866_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2866_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2866_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2866_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3037_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3037_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3037_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3037_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3037_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3049_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3049_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3049_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3049_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3049_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3322_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3322_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3322_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3322_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3322_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3322_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3406_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3406_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3406_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3406_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3406_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3430_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3430_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3430_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3430_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3430_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3430_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3624_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3624_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3624_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3624_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3624_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3636_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3636_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3636_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_3636_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3636_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3902_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3902_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3902_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3902_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3902_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3902_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3986_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3986_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3986_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3986_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3986_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4010_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4010_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4010_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4010_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4010_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4010_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4193_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4193_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4193_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4193_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4193_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4205_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4205_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4205_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4205_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4205_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4466_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4466_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4466_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4466_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4466_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4466_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4550_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4550_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4550_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4550_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4550_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4574_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_4574_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4574_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_4574_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_4574_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4574_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_4762_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4762_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4762_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4762_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4762_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4774_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_4774_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4774_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_4774_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_4774_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_5028_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_5028_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5028_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5028_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_5028_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5028_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5112_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_5112_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5112_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5112_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5112_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5136_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_5136_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5136_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_5136_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_5136_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_5136_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_727_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_727_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_727_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_727_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_727_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_746_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_746_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_746_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_746_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_746_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_765_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_765_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_765_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_765_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_765_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_794_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_794_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_794_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_794_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_794_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_806_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_806_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_806_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_806_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_806_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext1717_887 : std_logic_vector(31 downto 0);
    signal sext1718_1401 : std_logic_vector(31 downto 0);
    signal sext1719_1451 : std_logic_vector(31 downto 0);
    signal sext1720_1953 : std_logic_vector(31 downto 0);
    signal sext1721_2003 : std_logic_vector(31 downto 0);
    signal sext1722_2528 : std_logic_vector(31 downto 0);
    signal sext1723_2578 : std_logic_vector(31 downto 0);
    signal sext1724_3079 : std_logic_vector(31 downto 0);
    signal sext1725_3129 : std_logic_vector(31 downto 0);
    signal sext1726_3666 : std_logic_vector(31 downto 0);
    signal sext1727_3716 : std_logic_vector(31 downto 0);
    signal sext1728_4235 : std_logic_vector(31 downto 0);
    signal sext1729_4285 : std_logic_vector(31 downto 0);
    signal sext1730_4804 : std_logic_vector(31 downto 0);
    signal sext1731_4854 : std_logic_vector(31 downto 0);
    signal sext1764_821 : std_logic_vector(31 downto 0);
    signal sext1765_861 : std_logic_vector(31 downto 0);
    signal sext1766_1386 : std_logic_vector(31 downto 0);
    signal sext1767_1425 : std_logic_vector(31 downto 0);
    signal sext1768_1938 : std_logic_vector(31 downto 0);
    signal sext1769_1977 : std_logic_vector(31 downto 0);
    signal sext1770_2513 : std_logic_vector(31 downto 0);
    signal sext1771_2552 : std_logic_vector(31 downto 0);
    signal sext1772_3064 : std_logic_vector(31 downto 0);
    signal sext1773_3103 : std_logic_vector(31 downto 0);
    signal sext1774_3651 : std_logic_vector(31 downto 0);
    signal sext1775_3690 : std_logic_vector(31 downto 0);
    signal sext1776_4220 : std_logic_vector(31 downto 0);
    signal sext1777_4259 : std_logic_vector(31 downto 0);
    signal sext1778_4789 : std_logic_vector(31 downto 0);
    signal sext1779_4828 : std_logic_vector(31 downto 0);
    signal sext_837 : std_logic_vector(31 downto 0);
    signal shl1029_3118 : std_logic_vector(31 downto 0);
    signal shl1251_3705 : std_logic_vector(31 downto 0);
    signal shl1470_4274 : std_logic_vector(31 downto 0);
    signal shl1689_4843 : std_logic_vector(31 downto 0);
    signal shl372_1440 : std_logic_vector(31 downto 0);
    signal shl590_1992 : std_logic_vector(31 downto 0);
    signal shl810_2567 : std_logic_vector(31 downto 0);
    signal shl_876 : std_logic_vector(31 downto 0);
    signal shr1001_3416 : std_logic_vector(31 downto 0);
    signal shr1176_3888 : std_logic_vector(31 downto 0);
    signal shr1219_3971 : std_logic_vector(31 downto 0);
    signal shr1224_3996 : std_logic_vector(31 downto 0);
    signal shr129_1145 : std_logic_vector(31 downto 0);
    signal shr134_1170 : std_logic_vector(31 downto 0);
    signal shr1394_4452 : std_logic_vector(31 downto 0);
    signal shr1437_4535 : std_logic_vector(31 downto 0);
    signal shr1442_4560 : std_logic_vector(31 downto 0);
    signal shr1614_5014 : std_logic_vector(31 downto 0);
    signal shr1657_5097 : std_logic_vector(31 downto 0);
    signal shr1662_5122 : std_logic_vector(31 downto 0);
    signal shr297_1618 : std_logic_vector(31 downto 0);
    signal shr340_1701 : std_logic_vector(31 downto 0);
    signal shr345_1726 : std_logic_vector(31 downto 0);
    signal shr514_2176 : std_logic_vector(31 downto 0);
    signal shr557_2259 : std_logic_vector(31 downto 0);
    signal shr562_2284 : std_logic_vector(31 downto 0);
    signal shr735_2744 : std_logic_vector(31 downto 0);
    signal shr778_2827 : std_logic_vector(31 downto 0);
    signal shr783_2852 : std_logic_vector(31 downto 0);
    signal shr953_3308 : std_logic_vector(31 downto 0);
    signal shr996_3391 : std_logic_vector(31 downto 0);
    signal shr_1061 : std_logic_vector(31 downto 0);
    signal sub109_1101 : std_logic_vector(31 downto 0);
    signal sub1190_3917 : std_logic_vector(31 downto 0);
    signal sub1199_3927 : std_logic_vector(31 downto 0);
    signal sub1408_4481 : std_logic_vector(31 downto 0);
    signal sub1417_4491 : std_logic_vector(31 downto 0);
    signal sub1628_5043 : std_logic_vector(31 downto 0);
    signal sub1637_5053 : std_logic_vector(31 downto 0);
    signal sub311_1647 : std_logic_vector(31 downto 0);
    signal sub320_1657 : std_logic_vector(31 downto 0);
    signal sub528_2205 : std_logic_vector(31 downto 0);
    signal sub537_2215 : std_logic_vector(31 downto 0);
    signal sub749_2773 : std_logic_vector(31 downto 0);
    signal sub758_2783 : std_logic_vector(31 downto 0);
    signal sub967_3337 : std_logic_vector(31 downto 0);
    signal sub976_3347 : std_logic_vector(31 downto 0);
    signal sub_1091 : std_logic_vector(31 downto 0);
    signal tmp1024_3481 : std_logic_vector(7 downto 0);
    signal tmp1040_3525 : std_logic_vector(7 downto 0);
    signal tmp1063_3584 : std_logic_vector(7 downto 0);
    signal tmp1069_3597 : std_logic_vector(7 downto 0);
    signal tmp1075_3610 : std_logic_vector(7 downto 0);
    signal tmp1079_3613 : std_logic_vector(7 downto 0);
    signal tmp1091_3625 : std_logic_vector(31 downto 0);
    signal tmp1095_3637 : std_logic_vector(31 downto 0);
    signal tmp1132_3769 : std_logic_vector(7 downto 0);
    signal tmp1151_3826 : std_logic_vector(7 downto 0);
    signal tmp1222_3987 : std_logic_vector(63 downto 0);
    signal tmp1247_4061 : std_logic_vector(7 downto 0);
    signal tmp1262_4098 : std_logic_vector(7 downto 0);
    signal tmp1287_4157 : std_logic_vector(7 downto 0);
    signal tmp1294_4176 : std_logic_vector(7 downto 0);
    signal tmp1298_4179 : std_logic_vector(7 downto 0);
    signal tmp12_780 : std_logic_vector(7 downto 0);
    signal tmp1302_4182 : std_logic_vector(7 downto 0);
    signal tmp1310_4194 : std_logic_vector(31 downto 0);
    signal tmp1314_4206 : std_logic_vector(31 downto 0);
    signal tmp132_1161 : std_logic_vector(63 downto 0);
    signal tmp1351_4339 : std_logic_vector(7 downto 0);
    signal tmp1368_4384 : std_logic_vector(7 downto 0);
    signal tmp1440_4551 : std_logic_vector(63 downto 0);
    signal tmp1465_4625 : std_logic_vector(7 downto 0);
    signal tmp1481_4669 : std_logic_vector(7 downto 0);
    signal tmp1502_4716 : std_logic_vector(7 downto 0);
    signal tmp1508_4729 : std_logic_vector(7 downto 0);
    signal tmp1515_4748 : std_logic_vector(7 downto 0);
    signal tmp1519_4751 : std_logic_vector(7 downto 0);
    signal tmp1531_4763 : std_logic_vector(31 downto 0);
    signal tmp1535_4775 : std_logic_vector(31 downto 0);
    signal tmp154_1235 : std_logic_vector(7 downto 0);
    signal tmp1572_4907 : std_logic_vector(7 downto 0);
    signal tmp1589_4952 : std_logic_vector(7 downto 0);
    signal tmp15_783 : std_logic_vector(7 downto 0);
    signal tmp1660_5113 : std_logic_vector(63 downto 0);
    signal tmp1685_5187 : std_logic_vector(7 downto 0);
    signal tmp169_1279 : std_logic_vector(7 downto 0);
    signal tmp1700_5224 : std_logic_vector(7 downto 0);
    signal tmp189_1332 : std_logic_vector(7 downto 0);
    signal tmp197_1345 : std_logic_vector(7 downto 0);
    signal tmp1_747 : std_logic_vector(31 downto 0);
    signal tmp201_1348 : std_logic_vector(7 downto 0);
    signal tmp213_1360 : std_logic_vector(31 downto 0);
    signal tmp217_1372 : std_logic_vector(31 downto 0);
    signal tmp21_795 : std_logic_vector(31 downto 0);
    signal tmp24_807 : std_logic_vector(31 downto 0);
    signal tmp254_1505 : std_logic_vector(7 downto 0);
    signal tmp272_1556 : std_logic_vector(7 downto 0);
    signal tmp343_1717 : std_logic_vector(63 downto 0);
    signal tmp368_1791 : std_logic_vector(7 downto 0);
    signal tmp383_1828 : std_logic_vector(7 downto 0);
    signal tmp3_766 : std_logic_vector(31 downto 0);
    signal tmp407_1881 : std_logic_vector(7 downto 0);
    signal tmp413_1894 : std_logic_vector(7 downto 0);
    signal tmp417_1897 : std_logic_vector(7 downto 0);
    signal tmp421_1900 : std_logic_vector(7 downto 0);
    signal tmp429_1912 : std_logic_vector(31 downto 0);
    signal tmp433_1924 : std_logic_vector(31 downto 0);
    signal tmp470_2057 : std_logic_vector(7 downto 0);
    signal tmp488_2108 : std_logic_vector(7 downto 0);
    signal tmp52_942 : std_logic_vector(7 downto 0);
    signal tmp560_2275 : std_logic_vector(63 downto 0);
    signal tmp585_2349 : std_logic_vector(7 downto 0);
    signal tmp601_2393 : std_logic_vector(7 downto 0);
    signal tmp623_2446 : std_logic_vector(7 downto 0);
    signal tmp629_2459 : std_logic_vector(7 downto 0);
    signal tmp635_2472 : std_logic_vector(7 downto 0);
    signal tmp639_2475 : std_logic_vector(7 downto 0);
    signal tmp651_2487 : std_logic_vector(31 downto 0);
    signal tmp655_2499 : std_logic_vector(31 downto 0);
    signal tmp68_993 : std_logic_vector(7 downto 0);
    signal tmp692_2631 : std_logic_vector(7 downto 0);
    signal tmp710_2682 : std_logic_vector(7 downto 0);
    signal tmp781_2843 : std_logic_vector(63 downto 0);
    signal tmp806_2917 : std_logic_vector(7 downto 0);
    signal tmp821_2954 : std_logic_vector(7 downto 0);
    signal tmp845_3007 : std_logic_vector(7 downto 0);
    signal tmp851_3020 : std_logic_vector(7 downto 0);
    signal tmp855_3023 : std_logic_vector(7 downto 0);
    signal tmp859_3026 : std_logic_vector(7 downto 0);
    signal tmp867_3038 : std_logic_vector(31 downto 0);
    signal tmp871_3050 : std_logic_vector(31 downto 0);
    signal tmp908_3183 : std_logic_vector(7 downto 0);
    signal tmp927_3240 : std_logic_vector(7 downto 0);
    signal tmp999_3407 : std_logic_vector(63 downto 0);
    signal tmp9_777 : std_logic_vector(7 downto 0);
    signal tmp_728 : std_logic_vector(31 downto 0);
    signal type_cast_1001_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1011_wire : std_logic_vector(31 downto 0);
    signal type_cast_1013_wire : std_logic_vector(31 downto 0);
    signal type_cast_1025_wire : std_logic_vector(31 downto 0);
    signal type_cast_1030_wire : std_logic_vector(31 downto 0);
    signal type_cast_1055_wire : std_logic_vector(31 downto 0);
    signal type_cast_1058_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1065_wire : std_logic_vector(63 downto 0);
    signal type_cast_1078_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1084_wire : std_logic_vector(31 downto 0);
    signal type_cast_1139_wire : std_logic_vector(31 downto 0);
    signal type_cast_1142_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1148_wire : std_logic_vector(63 downto 0);
    signal type_cast_1164_wire : std_logic_vector(31 downto 0);
    signal type_cast_1167_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1173_wire : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire : std_logic_vector(31 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1202_wire : std_logic_vector(31 downto 0);
    signal type_cast_1204_wire : std_logic_vector(31 downto 0);
    signal type_cast_1217_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1230_wire : std_logic_vector(31 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1274_wire : std_logic_vector(31 downto 0);
    signal type_cast_1287_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1310_wire : std_logic_vector(15 downto 0);
    signal type_cast_1312_wire : std_logic_vector(15 downto 0);
    signal type_cast_1316_wire : std_logic_vector(15 downto 0);
    signal type_cast_1318_wire : std_logic_vector(15 downto 0);
    signal type_cast_1323_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1325_wire : std_logic_vector(15 downto 0);
    signal type_cast_1340_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1384_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1389_wire : std_logic_vector(31 downto 0);
    signal type_cast_1392_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1399_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1404_wire : std_logic_vector(31 downto 0);
    signal type_cast_1407_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1423_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1428_wire : std_logic_vector(31 downto 0);
    signal type_cast_1431_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1444_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1454_wire : std_logic_vector(31 downto 0);
    signal type_cast_1457_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1466_wire : std_logic_vector(15 downto 0);
    signal type_cast_1468_wire : std_logic_vector(15 downto 0);
    signal type_cast_1473_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1475_wire : std_logic_vector(15 downto 0);
    signal type_cast_1480_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1482_wire : std_logic_vector(15 downto 0);
    signal type_cast_1486_wire : std_logic_vector(31 downto 0);
    signal type_cast_1491_wire : std_logic_vector(31 downto 0);
    signal type_cast_1493_wire : std_logic_vector(31 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1523_wire : std_logic_vector(31 downto 0);
    signal type_cast_1525_wire : std_logic_vector(31 downto 0);
    signal type_cast_1537_wire : std_logic_vector(31 downto 0);
    signal type_cast_1542_wire : std_logic_vector(31 downto 0);
    signal type_cast_1544_wire : std_logic_vector(31 downto 0);
    signal type_cast_1568_wire : std_logic_vector(31 downto 0);
    signal type_cast_1570_wire : std_logic_vector(31 downto 0);
    signal type_cast_1582_wire : std_logic_vector(31 downto 0);
    signal type_cast_1587_wire : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire : std_logic_vector(31 downto 0);
    signal type_cast_1615_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1621_wire : std_logic_vector(63 downto 0);
    signal type_cast_1634_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1640_wire : std_logic_vector(31 downto 0);
    signal type_cast_1695_wire : std_logic_vector(31 downto 0);
    signal type_cast_1698_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1704_wire : std_logic_vector(63 downto 0);
    signal type_cast_1720_wire : std_logic_vector(31 downto 0);
    signal type_cast_1723_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1729_wire : std_logic_vector(63 downto 0);
    signal type_cast_1747_wire : std_logic_vector(31 downto 0);
    signal type_cast_1753_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1758_wire : std_logic_vector(31 downto 0);
    signal type_cast_1760_wire : std_logic_vector(31 downto 0);
    signal type_cast_1773_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1781_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1786_wire : std_logic_vector(31 downto 0);
    signal type_cast_1823_wire : std_logic_vector(31 downto 0);
    signal type_cast_1836_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1859_wire : std_logic_vector(15 downto 0);
    signal type_cast_1861_wire : std_logic_vector(15 downto 0);
    signal type_cast_1865_wire : std_logic_vector(15 downto 0);
    signal type_cast_1867_wire : std_logic_vector(15 downto 0);
    signal type_cast_1871_wire : std_logic_vector(15 downto 0);
    signal type_cast_1874_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1889_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1936_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1941_wire : std_logic_vector(31 downto 0);
    signal type_cast_1944_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1951_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1956_wire : std_logic_vector(31 downto 0);
    signal type_cast_1959_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1975_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1980_wire : std_logic_vector(31 downto 0);
    signal type_cast_1983_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1990_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1996_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2006_wire : std_logic_vector(31 downto 0);
    signal type_cast_2009_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2018_wire : std_logic_vector(15 downto 0);
    signal type_cast_2021_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2025_wire : std_logic_vector(15 downto 0);
    signal type_cast_2027_wire : std_logic_vector(15 downto 0);
    signal type_cast_2031_wire : std_logic_vector(15 downto 0);
    signal type_cast_2034_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2038_wire : std_logic_vector(31 downto 0);
    signal type_cast_2043_wire : std_logic_vector(31 downto 0);
    signal type_cast_2045_wire : std_logic_vector(31 downto 0);
    signal type_cast_2065_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2075_wire : std_logic_vector(31 downto 0);
    signal type_cast_2077_wire : std_logic_vector(31 downto 0);
    signal type_cast_2089_wire : std_logic_vector(31 downto 0);
    signal type_cast_2094_wire : std_logic_vector(31 downto 0);
    signal type_cast_2096_wire : std_logic_vector(31 downto 0);
    signal type_cast_2116_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2126_wire : std_logic_vector(31 downto 0);
    signal type_cast_2128_wire : std_logic_vector(31 downto 0);
    signal type_cast_2140_wire : std_logic_vector(31 downto 0);
    signal type_cast_2145_wire : std_logic_vector(31 downto 0);
    signal type_cast_2170_wire : std_logic_vector(31 downto 0);
    signal type_cast_2173_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2179_wire : std_logic_vector(63 downto 0);
    signal type_cast_2192_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2198_wire : std_logic_vector(31 downto 0);
    signal type_cast_2253_wire : std_logic_vector(31 downto 0);
    signal type_cast_2256_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2262_wire : std_logic_vector(63 downto 0);
    signal type_cast_2278_wire : std_logic_vector(31 downto 0);
    signal type_cast_2281_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2287_wire : std_logic_vector(63 downto 0);
    signal type_cast_2305_wire : std_logic_vector(31 downto 0);
    signal type_cast_2311_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2316_wire : std_logic_vector(31 downto 0);
    signal type_cast_2318_wire : std_logic_vector(31 downto 0);
    signal type_cast_2331_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2339_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2344_wire : std_logic_vector(31 downto 0);
    signal type_cast_2357_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2382_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2388_wire : std_logic_vector(31 downto 0);
    signal type_cast_2401_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2424_wire : std_logic_vector(15 downto 0);
    signal type_cast_2427_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2431_wire : std_logic_vector(15 downto 0);
    signal type_cast_2433_wire : std_logic_vector(15 downto 0);
    signal type_cast_2437_wire : std_logic_vector(15 downto 0);
    signal type_cast_2439_wire : std_logic_vector(15 downto 0);
    signal type_cast_2454_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2467_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2511_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2516_wire : std_logic_vector(31 downto 0);
    signal type_cast_2519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2526_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2531_wire : std_logic_vector(31 downto 0);
    signal type_cast_2534_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2550_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2555_wire : std_logic_vector(31 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2565_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2571_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2581_wire : std_logic_vector(31 downto 0);
    signal type_cast_2584_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2596_wire : std_logic_vector(15 downto 0);
    signal type_cast_2600_wire : std_logic_vector(15 downto 0);
    signal type_cast_2602_wire : std_logic_vector(15 downto 0);
    signal type_cast_2606_wire : std_logic_vector(15 downto 0);
    signal type_cast_2608_wire : std_logic_vector(15 downto 0);
    signal type_cast_2612_wire : std_logic_vector(31 downto 0);
    signal type_cast_2617_wire : std_logic_vector(31 downto 0);
    signal type_cast_2619_wire : std_logic_vector(31 downto 0);
    signal type_cast_2639_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2649_wire : std_logic_vector(31 downto 0);
    signal type_cast_2651_wire : std_logic_vector(31 downto 0);
    signal type_cast_2663_wire : std_logic_vector(31 downto 0);
    signal type_cast_2668_wire : std_logic_vector(31 downto 0);
    signal type_cast_2670_wire : std_logic_vector(31 downto 0);
    signal type_cast_2694_wire : std_logic_vector(31 downto 0);
    signal type_cast_2696_wire : std_logic_vector(31 downto 0);
    signal type_cast_2708_wire : std_logic_vector(31 downto 0);
    signal type_cast_2713_wire : std_logic_vector(31 downto 0);
    signal type_cast_2738_wire : std_logic_vector(31 downto 0);
    signal type_cast_2741_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2747_wire : std_logic_vector(63 downto 0);
    signal type_cast_2760_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2766_wire : std_logic_vector(31 downto 0);
    signal type_cast_2821_wire : std_logic_vector(31 downto 0);
    signal type_cast_2824_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2830_wire : std_logic_vector(63 downto 0);
    signal type_cast_2846_wire : std_logic_vector(31 downto 0);
    signal type_cast_2849_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2855_wire : std_logic_vector(63 downto 0);
    signal type_cast_2873_wire : std_logic_vector(31 downto 0);
    signal type_cast_2879_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2884_wire : std_logic_vector(31 downto 0);
    signal type_cast_2886_wire : std_logic_vector(31 downto 0);
    signal type_cast_2899_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2907_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2912_wire : std_logic_vector(31 downto 0);
    signal type_cast_2949_wire : std_logic_vector(31 downto 0);
    signal type_cast_2962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2985_wire : std_logic_vector(15 downto 0);
    signal type_cast_2988_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2992_wire : std_logic_vector(15 downto 0);
    signal type_cast_2994_wire : std_logic_vector(15 downto 0);
    signal type_cast_2998_wire : std_logic_vector(15 downto 0);
    signal type_cast_3000_wire : std_logic_vector(15 downto 0);
    signal type_cast_3015_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3062_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3067_wire : std_logic_vector(31 downto 0);
    signal type_cast_3070_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3077_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3082_wire : std_logic_vector(31 downto 0);
    signal type_cast_3085_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3101_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3106_wire : std_logic_vector(31 downto 0);
    signal type_cast_3109_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3116_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3122_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3132_wire : std_logic_vector(31 downto 0);
    signal type_cast_3135_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3144_wire : std_logic_vector(15 downto 0);
    signal type_cast_3147_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3151_wire : std_logic_vector(15 downto 0);
    signal type_cast_3153_wire : std_logic_vector(15 downto 0);
    signal type_cast_3157_wire : std_logic_vector(15 downto 0);
    signal type_cast_3160_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3164_wire : std_logic_vector(31 downto 0);
    signal type_cast_3169_wire : std_logic_vector(31 downto 0);
    signal type_cast_3171_wire : std_logic_vector(31 downto 0);
    signal type_cast_3191_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3207_wire : std_logic_vector(31 downto 0);
    signal type_cast_3209_wire : std_logic_vector(31 downto 0);
    signal type_cast_3221_wire : std_logic_vector(31 downto 0);
    signal type_cast_3226_wire : std_logic_vector(31 downto 0);
    signal type_cast_3228_wire : std_logic_vector(31 downto 0);
    signal type_cast_3248_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3258_wire : std_logic_vector(31 downto 0);
    signal type_cast_3260_wire : std_logic_vector(31 downto 0);
    signal type_cast_3272_wire : std_logic_vector(31 downto 0);
    signal type_cast_3277_wire : std_logic_vector(31 downto 0);
    signal type_cast_3302_wire : std_logic_vector(31 downto 0);
    signal type_cast_3305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3311_wire : std_logic_vector(63 downto 0);
    signal type_cast_3324_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3330_wire : std_logic_vector(31 downto 0);
    signal type_cast_3385_wire : std_logic_vector(31 downto 0);
    signal type_cast_3388_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3394_wire : std_logic_vector(63 downto 0);
    signal type_cast_3410_wire : std_logic_vector(31 downto 0);
    signal type_cast_3413_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3419_wire : std_logic_vector(63 downto 0);
    signal type_cast_3437_wire : std_logic_vector(31 downto 0);
    signal type_cast_3443_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3448_wire : std_logic_vector(31 downto 0);
    signal type_cast_3450_wire : std_logic_vector(31 downto 0);
    signal type_cast_3463_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3471_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3476_wire : std_logic_vector(31 downto 0);
    signal type_cast_3489_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3514_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3520_wire : std_logic_vector(31 downto 0);
    signal type_cast_3533_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3539_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3562_wire : std_logic_vector(15 downto 0);
    signal type_cast_3565_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3569_wire : std_logic_vector(15 downto 0);
    signal type_cast_3571_wire : std_logic_vector(15 downto 0);
    signal type_cast_3575_wire : std_logic_vector(15 downto 0);
    signal type_cast_3577_wire : std_logic_vector(15 downto 0);
    signal type_cast_3592_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3605_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3654_wire : std_logic_vector(31 downto 0);
    signal type_cast_3657_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3669_wire : std_logic_vector(31 downto 0);
    signal type_cast_3672_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3688_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3693_wire : std_logic_vector(31 downto 0);
    signal type_cast_3696_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3703_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3709_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3719_wire : std_logic_vector(31 downto 0);
    signal type_cast_3722_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3731_wire : std_logic_vector(15 downto 0);
    signal type_cast_3734_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3738_wire : std_logic_vector(15 downto 0);
    signal type_cast_3740_wire : std_logic_vector(15 downto 0);
    signal type_cast_3744_wire : std_logic_vector(15 downto 0);
    signal type_cast_3746_wire : std_logic_vector(15 downto 0);
    signal type_cast_3750_wire : std_logic_vector(31 downto 0);
    signal type_cast_3755_wire : std_logic_vector(31 downto 0);
    signal type_cast_3757_wire : std_logic_vector(31 downto 0);
    signal type_cast_3777_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3783_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3793_wire : std_logic_vector(31 downto 0);
    signal type_cast_3795_wire : std_logic_vector(31 downto 0);
    signal type_cast_3807_wire : std_logic_vector(31 downto 0);
    signal type_cast_3812_wire : std_logic_vector(31 downto 0);
    signal type_cast_3814_wire : std_logic_vector(31 downto 0);
    signal type_cast_3838_wire : std_logic_vector(31 downto 0);
    signal type_cast_3840_wire : std_logic_vector(31 downto 0);
    signal type_cast_3852_wire : std_logic_vector(31 downto 0);
    signal type_cast_3857_wire : std_logic_vector(31 downto 0);
    signal type_cast_3882_wire : std_logic_vector(31 downto 0);
    signal type_cast_3885_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3891_wire : std_logic_vector(63 downto 0);
    signal type_cast_3904_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3910_wire : std_logic_vector(31 downto 0);
    signal type_cast_3965_wire : std_logic_vector(31 downto 0);
    signal type_cast_3968_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3974_wire : std_logic_vector(63 downto 0);
    signal type_cast_3990_wire : std_logic_vector(31 downto 0);
    signal type_cast_3993_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3999_wire : std_logic_vector(63 downto 0);
    signal type_cast_4017_wire : std_logic_vector(31 downto 0);
    signal type_cast_4023_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4028_wire : std_logic_vector(31 downto 0);
    signal type_cast_4030_wire : std_logic_vector(31 downto 0);
    signal type_cast_4043_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4051_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4056_wire : std_logic_vector(31 downto 0);
    signal type_cast_4093_wire : std_logic_vector(31 downto 0);
    signal type_cast_4106_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4112_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4135_wire : std_logic_vector(15 downto 0);
    signal type_cast_4138_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4142_wire : std_logic_vector(15 downto 0);
    signal type_cast_4144_wire : std_logic_vector(15 downto 0);
    signal type_cast_4148_wire : std_logic_vector(15 downto 0);
    signal type_cast_4150_wire : std_logic_vector(15 downto 0);
    signal type_cast_4165_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4171_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4218_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4223_wire : std_logic_vector(31 downto 0);
    signal type_cast_4226_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4238_wire : std_logic_vector(31 downto 0);
    signal type_cast_4241_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4257_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4262_wire : std_logic_vector(31 downto 0);
    signal type_cast_4265_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4272_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4278_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4288_wire : std_logic_vector(31 downto 0);
    signal type_cast_4291_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4301_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4303_wire : std_logic_vector(15 downto 0);
    signal type_cast_4307_wire : std_logic_vector(15 downto 0);
    signal type_cast_4309_wire : std_logic_vector(15 downto 0);
    signal type_cast_4314_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4316_wire : std_logic_vector(15 downto 0);
    signal type_cast_4320_wire : std_logic_vector(31 downto 0);
    signal type_cast_4325_wire : std_logic_vector(31 downto 0);
    signal type_cast_4327_wire : std_logic_vector(31 downto 0);
    signal type_cast_4351_wire : std_logic_vector(31 downto 0);
    signal type_cast_4353_wire : std_logic_vector(31 downto 0);
    signal type_cast_4365_wire : std_logic_vector(31 downto 0);
    signal type_cast_4370_wire : std_logic_vector(31 downto 0);
    signal type_cast_4372_wire : std_logic_vector(31 downto 0);
    signal type_cast_4392_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4402_wire : std_logic_vector(31 downto 0);
    signal type_cast_4404_wire : std_logic_vector(31 downto 0);
    signal type_cast_4416_wire : std_logic_vector(31 downto 0);
    signal type_cast_4421_wire : std_logic_vector(31 downto 0);
    signal type_cast_4446_wire : std_logic_vector(31 downto 0);
    signal type_cast_4449_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4455_wire : std_logic_vector(63 downto 0);
    signal type_cast_4468_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_4474_wire : std_logic_vector(31 downto 0);
    signal type_cast_4529_wire : std_logic_vector(31 downto 0);
    signal type_cast_4532_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4538_wire : std_logic_vector(63 downto 0);
    signal type_cast_4554_wire : std_logic_vector(31 downto 0);
    signal type_cast_4557_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4563_wire : std_logic_vector(63 downto 0);
    signal type_cast_4581_wire : std_logic_vector(31 downto 0);
    signal type_cast_4587_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4592_wire : std_logic_vector(31 downto 0);
    signal type_cast_4594_wire : std_logic_vector(31 downto 0);
    signal type_cast_4607_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4615_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4620_wire : std_logic_vector(31 downto 0);
    signal type_cast_4633_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4658_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4664_wire : std_logic_vector(31 downto 0);
    signal type_cast_4694_wire : std_logic_vector(15 downto 0);
    signal type_cast_4697_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4701_wire : std_logic_vector(15 downto 0);
    signal type_cast_4703_wire : std_logic_vector(15 downto 0);
    signal type_cast_4707_wire : std_logic_vector(15 downto 0);
    signal type_cast_4709_wire : std_logic_vector(15 downto 0);
    signal type_cast_4724_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4737_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4743_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4787_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4792_wire : std_logic_vector(31 downto 0);
    signal type_cast_4795_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4802_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4807_wire : std_logic_vector(31 downto 0);
    signal type_cast_4810_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4826_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4831_wire : std_logic_vector(31 downto 0);
    signal type_cast_4834_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4841_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4847_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4857_wire : std_logic_vector(31 downto 0);
    signal type_cast_4860_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_4870_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_4872_wire : std_logic_vector(15 downto 0);
    signal type_cast_4876_wire : std_logic_vector(15 downto 0);
    signal type_cast_4878_wire : std_logic_vector(15 downto 0);
    signal type_cast_4882_wire : std_logic_vector(15 downto 0);
    signal type_cast_4884_wire : std_logic_vector(15 downto 0);
    signal type_cast_4888_wire : std_logic_vector(31 downto 0);
    signal type_cast_4893_wire : std_logic_vector(31 downto 0);
    signal type_cast_4895_wire : std_logic_vector(31 downto 0);
    signal type_cast_4919_wire : std_logic_vector(31 downto 0);
    signal type_cast_4921_wire : std_logic_vector(31 downto 0);
    signal type_cast_4933_wire : std_logic_vector(31 downto 0);
    signal type_cast_4938_wire : std_logic_vector(31 downto 0);
    signal type_cast_4940_wire : std_logic_vector(31 downto 0);
    signal type_cast_4964_wire : std_logic_vector(31 downto 0);
    signal type_cast_4966_wire : std_logic_vector(31 downto 0);
    signal type_cast_4978_wire : std_logic_vector(31 downto 0);
    signal type_cast_4983_wire : std_logic_vector(31 downto 0);
    signal type_cast_5008_wire : std_logic_vector(31 downto 0);
    signal type_cast_5011_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5017_wire : std_logic_vector(63 downto 0);
    signal type_cast_5030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_5036_wire : std_logic_vector(31 downto 0);
    signal type_cast_5091_wire : std_logic_vector(31 downto 0);
    signal type_cast_5094_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5100_wire : std_logic_vector(63 downto 0);
    signal type_cast_5116_wire : std_logic_vector(31 downto 0);
    signal type_cast_5119_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5125_wire : std_logic_vector(63 downto 0);
    signal type_cast_5143_wire : std_logic_vector(31 downto 0);
    signal type_cast_5149_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_5154_wire : std_logic_vector(31 downto 0);
    signal type_cast_5156_wire : std_logic_vector(31 downto 0);
    signal type_cast_5169_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_5177_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_5182_wire : std_logic_vector(31 downto 0);
    signal type_cast_5219_wire : std_logic_vector(31 downto 0);
    signal type_cast_5250_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_5252_wire : std_logic_vector(15 downto 0);
    signal type_cast_5256_wire : std_logic_vector(15 downto 0);
    signal type_cast_5258_wire : std_logic_vector(15 downto 0);
    signal type_cast_5262_wire : std_logic_vector(15 downto 0);
    signal type_cast_5264_wire : std_logic_vector(15 downto 0);
    signal type_cast_819_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_825_wire : std_logic_vector(31 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_840_wire : std_logic_vector(31 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_864_wire : std_logic_vector(31 downto 0);
    signal type_cast_867_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_880_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_890_wire : std_logic_vector(31 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_905_wire : std_logic_vector(15 downto 0);
    signal type_cast_910_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_912_wire : std_logic_vector(15 downto 0);
    signal type_cast_917_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_919_wire : std_logic_vector(15 downto 0);
    signal type_cast_923_wire : std_logic_vector(31 downto 0);
    signal type_cast_928_wire : std_logic_vector(31 downto 0);
    signal type_cast_930_wire : std_logic_vector(31 downto 0);
    signal type_cast_950_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_960_wire : std_logic_vector(31 downto 0);
    signal type_cast_962_wire : std_logic_vector(31 downto 0);
    signal type_cast_974_wire : std_logic_vector(31 downto 0);
    signal type_cast_979_wire : std_logic_vector(31 downto 0);
    signal type_cast_981_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_col_high_1234_word_address_0 <= "0";
    LOAD_col_high_1331_word_address_0 <= "0";
    LOAD_col_high_1555_word_address_0 <= "0";
    LOAD_col_high_1790_word_address_0 <= "0";
    LOAD_col_high_1899_word_address_0 <= "0";
    LOAD_col_high_2107_word_address_0 <= "0";
    LOAD_col_high_2348_word_address_0 <= "0";
    LOAD_col_high_2445_word_address_0 <= "0";
    LOAD_col_high_2681_word_address_0 <= "0";
    LOAD_col_high_2916_word_address_0 <= "0";
    LOAD_col_high_3025_word_address_0 <= "0";
    LOAD_col_high_3239_word_address_0 <= "0";
    LOAD_col_high_3480_word_address_0 <= "0";
    LOAD_col_high_3583_word_address_0 <= "0";
    LOAD_col_high_3825_word_address_0 <= "0";
    LOAD_col_high_4060_word_address_0 <= "0";
    LOAD_col_high_4181_word_address_0 <= "0";
    LOAD_col_high_4383_word_address_0 <= "0";
    LOAD_col_high_4624_word_address_0 <= "0";
    LOAD_col_high_4715_word_address_0 <= "0";
    LOAD_col_high_4951_word_address_0 <= "0";
    LOAD_col_high_5186_word_address_0 <= "0";
    LOAD_col_high_782_word_address_0 <= "0";
    LOAD_col_high_992_word_address_0 <= "0";
    LOAD_depth_high_1347_word_address_0 <= "0";
    LOAD_depth_high_1896_word_address_0 <= "0";
    LOAD_depth_high_2474_word_address_0 <= "0";
    LOAD_depth_high_3022_word_address_0 <= "0";
    LOAD_depth_high_3612_word_address_0 <= "0";
    LOAD_depth_high_4178_word_address_0 <= "0";
    LOAD_depth_high_4750_word_address_0 <= "0";
    LOAD_depth_high_779_word_address_0 <= "0";
    LOAD_pad_1344_word_address_0 <= "0";
    LOAD_pad_1893_word_address_0 <= "0";
    LOAD_pad_2471_word_address_0 <= "0";
    LOAD_pad_3019_word_address_0 <= "0";
    LOAD_pad_3609_word_address_0 <= "0";
    LOAD_pad_4175_word_address_0 <= "0";
    LOAD_pad_4747_word_address_0 <= "0";
    LOAD_pad_776_word_address_0 <= "0";
    LOAD_row_high_1278_word_address_0 <= "0";
    LOAD_row_high_1504_word_address_0 <= "0";
    LOAD_row_high_1827_word_address_0 <= "0";
    LOAD_row_high_1880_word_address_0 <= "0";
    LOAD_row_high_2056_word_address_0 <= "0";
    LOAD_row_high_2392_word_address_0 <= "0";
    LOAD_row_high_2458_word_address_0 <= "0";
    LOAD_row_high_2630_word_address_0 <= "0";
    LOAD_row_high_2953_word_address_0 <= "0";
    LOAD_row_high_3006_word_address_0 <= "0";
    LOAD_row_high_3182_word_address_0 <= "0";
    LOAD_row_high_3524_word_address_0 <= "0";
    LOAD_row_high_3596_word_address_0 <= "0";
    LOAD_row_high_3768_word_address_0 <= "0";
    LOAD_row_high_4097_word_address_0 <= "0";
    LOAD_row_high_4156_word_address_0 <= "0";
    LOAD_row_high_4338_word_address_0 <= "0";
    LOAD_row_high_4668_word_address_0 <= "0";
    LOAD_row_high_4728_word_address_0 <= "0";
    LOAD_row_high_4906_word_address_0 <= "0";
    LOAD_row_high_5223_word_address_0 <= "0";
    LOAD_row_high_941_word_address_0 <= "0";
    STORE_col_high_752_word_address_0 <= "0";
    STORE_depth_high_771_word_address_0 <= "0";
    STORE_row_high_733_word_address_0 <= "0";
    array_obj_ref_1072_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1072_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1072_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1072_resized_base_address <= "00000000000000";
    array_obj_ref_1155_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1155_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1155_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1155_resized_base_address <= "00000000000000";
    array_obj_ref_1180_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1180_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1180_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1180_resized_base_address <= "00000000000000";
    array_obj_ref_1628_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1628_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1628_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1628_resized_base_address <= "00000000000000";
    array_obj_ref_1711_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1711_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1711_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1711_resized_base_address <= "00000000000000";
    array_obj_ref_1736_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1736_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1736_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1736_resized_base_address <= "00000000000000";
    array_obj_ref_2186_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2186_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2186_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2186_resized_base_address <= "00000000000000";
    array_obj_ref_2269_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2269_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2269_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2269_resized_base_address <= "00000000000000";
    array_obj_ref_2294_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2294_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2294_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2294_resized_base_address <= "00000000000000";
    array_obj_ref_2754_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2754_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2754_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2754_resized_base_address <= "00000000000000";
    array_obj_ref_2837_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2837_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2837_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2837_resized_base_address <= "00000000000000";
    array_obj_ref_2862_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2862_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2862_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2862_resized_base_address <= "00000000000000";
    array_obj_ref_3318_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3318_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3318_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3318_resized_base_address <= "00000000000000";
    array_obj_ref_3401_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3401_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3401_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3401_resized_base_address <= "00000000000000";
    array_obj_ref_3426_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3426_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3426_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3426_resized_base_address <= "00000000000000";
    array_obj_ref_3898_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3898_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3898_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3898_resized_base_address <= "00000000000000";
    array_obj_ref_3981_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3981_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3981_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3981_resized_base_address <= "00000000000000";
    array_obj_ref_4006_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4006_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4006_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4006_resized_base_address <= "00000000000000";
    array_obj_ref_4462_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4462_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4462_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4462_resized_base_address <= "00000000000000";
    array_obj_ref_4545_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4545_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4545_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4545_resized_base_address <= "00000000000000";
    array_obj_ref_4570_constant_part_of_offset <= "00000000000000";
    array_obj_ref_4570_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_4570_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_4570_resized_base_address <= "00000000000000";
    array_obj_ref_5024_constant_part_of_offset <= "00000000000000";
    array_obj_ref_5024_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_5024_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_5024_resized_base_address <= "00000000000000";
    array_obj_ref_5107_constant_part_of_offset <= "00000000000000";
    array_obj_ref_5107_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_5107_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_5107_resized_base_address <= "00000000000000";
    array_obj_ref_5132_constant_part_of_offset <= "00000000000000";
    array_obj_ref_5132_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_5132_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_5132_resized_base_address <= "00000000000000";
    iNsTr_0_724 <= "00000000000000000000000000000011";
    iNsTr_107_4190 <= "00000000000000000000000000000101";
    iNsTr_108_4202 <= "00000000000000000000000000000100";
    iNsTr_124_4759 <= "00000000000000000000000000000101";
    iNsTr_125_4771 <= "00000000000000000000000000000100";
    iNsTr_22_1356 <= "00000000000000000000000000000101";
    iNsTr_23_1368 <= "00000000000000000000000000000100";
    iNsTr_2_743 <= "00000000000000000000000000000100";
    iNsTr_39_1908 <= "00000000000000000000000000000101";
    iNsTr_40_1920 <= "00000000000000000000000000000100";
    iNsTr_4_762 <= "00000000000000000000000000000101";
    iNsTr_56_2483 <= "00000000000000000000000000000101";
    iNsTr_57_2495 <= "00000000000000000000000000000100";
    iNsTr_73_3034 <= "00000000000000000000000000000101";
    iNsTr_74_3046 <= "00000000000000000000000000000100";
    iNsTr_7_791 <= "00000000000000000000000000000101";
    iNsTr_8_803 <= "00000000000000000000000000000100";
    iNsTr_90_3621 <= "00000000000000000000000000000101";
    iNsTr_91_3633 <= "00000000000000000000000000000100";
    ptr_deref_1076_word_offset_0 <= "00000000000000";
    ptr_deref_1160_word_offset_0 <= "00000000000000";
    ptr_deref_1184_word_offset_0 <= "00000000000000";
    ptr_deref_1359_word_offset_0 <= "0000000";
    ptr_deref_1371_word_offset_0 <= "0000000";
    ptr_deref_1632_word_offset_0 <= "00000000000000";
    ptr_deref_1716_word_offset_0 <= "00000000000000";
    ptr_deref_1740_word_offset_0 <= "00000000000000";
    ptr_deref_1911_word_offset_0 <= "0000000";
    ptr_deref_1923_word_offset_0 <= "0000000";
    ptr_deref_2190_word_offset_0 <= "00000000000000";
    ptr_deref_2274_word_offset_0 <= "00000000000000";
    ptr_deref_2298_word_offset_0 <= "00000000000000";
    ptr_deref_2486_word_offset_0 <= "0000000";
    ptr_deref_2498_word_offset_0 <= "0000000";
    ptr_deref_2758_word_offset_0 <= "00000000000000";
    ptr_deref_2842_word_offset_0 <= "00000000000000";
    ptr_deref_2866_word_offset_0 <= "00000000000000";
    ptr_deref_3037_word_offset_0 <= "0000000";
    ptr_deref_3049_word_offset_0 <= "0000000";
    ptr_deref_3322_word_offset_0 <= "00000000000000";
    ptr_deref_3406_word_offset_0 <= "00000000000000";
    ptr_deref_3430_word_offset_0 <= "00000000000000";
    ptr_deref_3624_word_offset_0 <= "0000000";
    ptr_deref_3636_word_offset_0 <= "0000000";
    ptr_deref_3902_word_offset_0 <= "00000000000000";
    ptr_deref_3986_word_offset_0 <= "00000000000000";
    ptr_deref_4010_word_offset_0 <= "00000000000000";
    ptr_deref_4193_word_offset_0 <= "0000000";
    ptr_deref_4205_word_offset_0 <= "0000000";
    ptr_deref_4466_word_offset_0 <= "00000000000000";
    ptr_deref_4550_word_offset_0 <= "00000000000000";
    ptr_deref_4574_word_offset_0 <= "00000000000000";
    ptr_deref_4762_word_offset_0 <= "0000000";
    ptr_deref_4774_word_offset_0 <= "0000000";
    ptr_deref_5028_word_offset_0 <= "00000000000000";
    ptr_deref_5112_word_offset_0 <= "00000000000000";
    ptr_deref_5136_word_offset_0 <= "00000000000000";
    ptr_deref_727_word_offset_0 <= "0000000";
    ptr_deref_746_word_offset_0 <= "0000000";
    ptr_deref_765_word_offset_0 <= "0000000";
    ptr_deref_794_word_offset_0 <= "0000000";
    ptr_deref_806_word_offset_0 <= "0000000";
    type_cast_1001_wire_constant <= "00000000000000000000000000000001";
    type_cast_1058_wire_constant <= "00000000000000000000000000000010";
    type_cast_1078_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1142_wire_constant <= "00000000000000000000000000000010";
    type_cast_1167_wire_constant <= "00000000000000000000000000000010";
    type_cast_1197_wire_constant <= "00000000000000000000000000000100";
    type_cast_1217_wire_constant <= "0000000000000100";
    type_cast_1225_wire_constant <= "0000000000000001";
    type_cast_1243_wire_constant <= "00000000000000000000000000000001";
    type_cast_1268_wire_constant <= "0000000000000000";
    type_cast_1287_wire_constant <= "00000000000000000000000000000010";
    type_cast_1323_wire_constant <= "0000000000000000";
    type_cast_1340_wire_constant <= "0000000000000001";
    type_cast_1384_wire_constant <= "00000000000000000000000000010000";
    type_cast_1392_wire_constant <= "00000000000000000000000000010000";
    type_cast_1399_wire_constant <= "00000000000000000000000000010000";
    type_cast_1407_wire_constant <= "00000000000000000000000000010000";
    type_cast_1423_wire_constant <= "00000000000000000000000000010000";
    type_cast_1431_wire_constant <= "00000000000000000000000000010000";
    type_cast_1438_wire_constant <= "00000000000000000000000000000001";
    type_cast_1444_wire_constant <= "00000000000000000000000000010000";
    type_cast_1457_wire_constant <= "00000000000000000000000000010000";
    type_cast_1473_wire_constant <= "0000000000000000";
    type_cast_1480_wire_constant <= "0000000000000000";
    type_cast_1513_wire_constant <= "00000000000000000000000000000010";
    type_cast_1615_wire_constant <= "00000000000000000000000000000010";
    type_cast_1634_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1698_wire_constant <= "00000000000000000000000000000010";
    type_cast_1723_wire_constant <= "00000000000000000000000000000010";
    type_cast_1753_wire_constant <= "00000000000000000000000000000100";
    type_cast_1773_wire_constant <= "0000000000000100";
    type_cast_1781_wire_constant <= "0000000000000001";
    type_cast_1836_wire_constant <= "00000000000000000000000000000010";
    type_cast_1874_wire_constant <= "0000000000000000";
    type_cast_1889_wire_constant <= "0000000000000010";
    type_cast_1936_wire_constant <= "00000000000000000000000000010000";
    type_cast_1944_wire_constant <= "00000000000000000000000000010000";
    type_cast_1951_wire_constant <= "00000000000000000000000000010000";
    type_cast_1959_wire_constant <= "00000000000000000000000000010000";
    type_cast_1975_wire_constant <= "00000000000000000000000000010000";
    type_cast_1983_wire_constant <= "00000000000000000000000000010000";
    type_cast_1990_wire_constant <= "00000000000000000000000000000001";
    type_cast_1996_wire_constant <= "00000000000000000000000000010000";
    type_cast_2009_wire_constant <= "00000000000000000000000000010000";
    type_cast_2021_wire_constant <= "0000000000000000";
    type_cast_2034_wire_constant <= "0000000000000000";
    type_cast_2065_wire_constant <= "00000000000000000000000000000001";
    type_cast_2116_wire_constant <= "00000000000000000000000000000001";
    type_cast_2173_wire_constant <= "00000000000000000000000000000010";
    type_cast_2192_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2256_wire_constant <= "00000000000000000000000000000010";
    type_cast_2281_wire_constant <= "00000000000000000000000000000010";
    type_cast_2311_wire_constant <= "00000000000000000000000000000100";
    type_cast_2331_wire_constant <= "0000000000000100";
    type_cast_2339_wire_constant <= "0000000000000001";
    type_cast_2357_wire_constant <= "00000000000000000000000000000001";
    type_cast_2382_wire_constant <= "0000000000000000";
    type_cast_2401_wire_constant <= "00000000000000000000000000000001";
    type_cast_2427_wire_constant <= "0000000000000000";
    type_cast_2454_wire_constant <= "0000000000000001";
    type_cast_2467_wire_constant <= "0000000000000010";
    type_cast_2511_wire_constant <= "00000000000000000000000000010000";
    type_cast_2519_wire_constant <= "00000000000000000000000000010000";
    type_cast_2526_wire_constant <= "00000000000000000000000000010000";
    type_cast_2534_wire_constant <= "00000000000000000000000000010000";
    type_cast_2550_wire_constant <= "00000000000000000000000000010000";
    type_cast_2558_wire_constant <= "00000000000000000000000000010000";
    type_cast_2565_wire_constant <= "00000000000000000000000000000001";
    type_cast_2571_wire_constant <= "00000000000000000000000000010000";
    type_cast_2584_wire_constant <= "00000000000000000000000000010000";
    type_cast_2594_wire_constant <= "0000000000000000";
    type_cast_2639_wire_constant <= "00000000000000000000000000000001";
    type_cast_2741_wire_constant <= "00000000000000000000000000000010";
    type_cast_2760_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2824_wire_constant <= "00000000000000000000000000000010";
    type_cast_2849_wire_constant <= "00000000000000000000000000000010";
    type_cast_2879_wire_constant <= "00000000000000000000000000000100";
    type_cast_2899_wire_constant <= "0000000000000100";
    type_cast_2907_wire_constant <= "0000000000000001";
    type_cast_2962_wire_constant <= "00000000000000000000000000000001";
    type_cast_2988_wire_constant <= "0000000000000000";
    type_cast_3015_wire_constant <= "0000000000000001";
    type_cast_3062_wire_constant <= "00000000000000000000000000010000";
    type_cast_3070_wire_constant <= "00000000000000000000000000010000";
    type_cast_3077_wire_constant <= "00000000000000000000000000010000";
    type_cast_3085_wire_constant <= "00000000000000000000000000010000";
    type_cast_3101_wire_constant <= "00000000000000000000000000010000";
    type_cast_3109_wire_constant <= "00000000000000000000000000010000";
    type_cast_3116_wire_constant <= "00000000000000000000000000000001";
    type_cast_3122_wire_constant <= "00000000000000000000000000010000";
    type_cast_3135_wire_constant <= "00000000000000000000000000010000";
    type_cast_3147_wire_constant <= "0000000000000000";
    type_cast_3160_wire_constant <= "0000000000000000";
    type_cast_3191_wire_constant <= "00000000000000000000000000000011";
    type_cast_3197_wire_constant <= "00000000000000000000000000000010";
    type_cast_3248_wire_constant <= "00000000000000000000000000000001";
    type_cast_3305_wire_constant <= "00000000000000000000000000000010";
    type_cast_3324_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3388_wire_constant <= "00000000000000000000000000000010";
    type_cast_3413_wire_constant <= "00000000000000000000000000000010";
    type_cast_3443_wire_constant <= "00000000000000000000000000000100";
    type_cast_3463_wire_constant <= "0000000000000100";
    type_cast_3471_wire_constant <= "0000000000000001";
    type_cast_3489_wire_constant <= "00000000000000000000000000000001";
    type_cast_3514_wire_constant <= "0000000000000000";
    type_cast_3533_wire_constant <= "00000000000000000000000000000011";
    type_cast_3539_wire_constant <= "00000000000000000000000000000010";
    type_cast_3565_wire_constant <= "0000000000000000";
    type_cast_3592_wire_constant <= "0000000000000001";
    type_cast_3605_wire_constant <= "0000000000000001";
    type_cast_3649_wire_constant <= "00000000000000000000000000010000";
    type_cast_3657_wire_constant <= "00000000000000000000000000010000";
    type_cast_3664_wire_constant <= "00000000000000000000000000010000";
    type_cast_3672_wire_constant <= "00000000000000000000000000010000";
    type_cast_3688_wire_constant <= "00000000000000000000000000010000";
    type_cast_3696_wire_constant <= "00000000000000000000000000010000";
    type_cast_3703_wire_constant <= "00000000000000000000000000000001";
    type_cast_3709_wire_constant <= "00000000000000000000000000010000";
    type_cast_3722_wire_constant <= "00000000000000000000000000010000";
    type_cast_3734_wire_constant <= "0000000000000000";
    type_cast_3777_wire_constant <= "00000000000000000000000000000011";
    type_cast_3783_wire_constant <= "00000000000000000000000000000010";
    type_cast_3885_wire_constant <= "00000000000000000000000000000010";
    type_cast_3904_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3968_wire_constant <= "00000000000000000000000000000010";
    type_cast_3993_wire_constant <= "00000000000000000000000000000010";
    type_cast_4023_wire_constant <= "00000000000000000000000000000100";
    type_cast_4043_wire_constant <= "0000000000000100";
    type_cast_4051_wire_constant <= "0000000000000001";
    type_cast_4106_wire_constant <= "00000000000000000000000000000011";
    type_cast_4112_wire_constant <= "00000000000000000000000000000010";
    type_cast_4138_wire_constant <= "0000000000000000";
    type_cast_4165_wire_constant <= "0000000000000010";
    type_cast_4171_wire_constant <= "0000000000000011";
    type_cast_4218_wire_constant <= "00000000000000000000000000010000";
    type_cast_4226_wire_constant <= "00000000000000000000000000010000";
    type_cast_4233_wire_constant <= "00000000000000000000000000010000";
    type_cast_4241_wire_constant <= "00000000000000000000000000010000";
    type_cast_4257_wire_constant <= "00000000000000000000000000010000";
    type_cast_4265_wire_constant <= "00000000000000000000000000010000";
    type_cast_4272_wire_constant <= "00000000000000000000000000000001";
    type_cast_4278_wire_constant <= "00000000000000000000000000010000";
    type_cast_4291_wire_constant <= "00000000000000000000000000010000";
    type_cast_4301_wire_constant <= "0000000000000000";
    type_cast_4314_wire_constant <= "0000000000000000";
    type_cast_4392_wire_constant <= "00000000000000000000000000000001";
    type_cast_4449_wire_constant <= "00000000000000000000000000000010";
    type_cast_4468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4532_wire_constant <= "00000000000000000000000000000010";
    type_cast_4557_wire_constant <= "00000000000000000000000000000010";
    type_cast_4587_wire_constant <= "00000000000000000000000000000100";
    type_cast_4607_wire_constant <= "0000000000000100";
    type_cast_4615_wire_constant <= "0000000000000001";
    type_cast_4633_wire_constant <= "00000000000000000000000000000001";
    type_cast_4658_wire_constant <= "0000000000000000";
    type_cast_4697_wire_constant <= "0000000000000000";
    type_cast_4724_wire_constant <= "0000000000000001";
    type_cast_4737_wire_constant <= "0000000000000011";
    type_cast_4743_wire_constant <= "0000000000000010";
    type_cast_4787_wire_constant <= "00000000000000000000000000010000";
    type_cast_4795_wire_constant <= "00000000000000000000000000010000";
    type_cast_4802_wire_constant <= "00000000000000000000000000010000";
    type_cast_4810_wire_constant <= "00000000000000000000000000010000";
    type_cast_4826_wire_constant <= "00000000000000000000000000010000";
    type_cast_4834_wire_constant <= "00000000000000000000000000010000";
    type_cast_4841_wire_constant <= "00000000000000000000000000000001";
    type_cast_4847_wire_constant <= "00000000000000000000000000010000";
    type_cast_4860_wire_constant <= "00000000000000000000000000010000";
    type_cast_4870_wire_constant <= "0000000000000000";
    type_cast_5011_wire_constant <= "00000000000000000000000000000010";
    type_cast_5030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_5094_wire_constant <= "00000000000000000000000000000010";
    type_cast_5119_wire_constant <= "00000000000000000000000000000010";
    type_cast_5149_wire_constant <= "00000000000000000000000000000100";
    type_cast_5169_wire_constant <= "0000000000000100";
    type_cast_5177_wire_constant <= "0000000000000001";
    type_cast_5250_wire_constant <= "0000000000000000";
    type_cast_819_wire_constant <= "00000000000000000000000000010000";
    type_cast_828_wire_constant <= "00000000000000000000000000010000";
    type_cast_835_wire_constant <= "00000000000000000000000000010000";
    type_cast_843_wire_constant <= "00000000000000000000000000010000";
    type_cast_859_wire_constant <= "00000000000000000000000000010000";
    type_cast_867_wire_constant <= "00000000000000000000000000010000";
    type_cast_874_wire_constant <= "00000000000000000000000000000001";
    type_cast_880_wire_constant <= "00000000000000000000000000010000";
    type_cast_893_wire_constant <= "00000000000000000000000000010000";
    type_cast_903_wire_constant <= "0000000000000000";
    type_cast_910_wire_constant <= "0000000000000000";
    type_cast_917_wire_constant <= "0000000000000000";
    type_cast_950_wire_constant <= "00000000000000000000000000000010";
    phi_stmt_1307: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1310_wire & type_cast_1312_wire;
      req <= phi_stmt_1307_req_0 & phi_stmt_1307_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1307",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1307_ack_0,
          idata => idata,
          odata => jx_x0x_xph_1307,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1307
    phi_stmt_1313: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1316_wire & type_cast_1318_wire;
      req <= phi_stmt_1313_req_0 & phi_stmt_1313_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1313",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1313_ack_0,
          idata => idata,
          odata => ix_x1x_xph_1313,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1313
    phi_stmt_1319: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1323_wire_constant & type_cast_1325_wire;
      req <= phi_stmt_1319_req_0 & phi_stmt_1319_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1319",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1319_ack_0,
          idata => idata,
          odata => kx_x0x_xph_1319,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1319
    phi_stmt_1463: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1466_wire & type_cast_1468_wire;
      req <= phi_stmt_1463_req_0 & phi_stmt_1463_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1463",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1463_ack_0,
          idata => idata,
          odata => j240x_x1_1463,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1463
    phi_stmt_1469: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1473_wire_constant & type_cast_1475_wire;
      req <= phi_stmt_1469_req_0 & phi_stmt_1469_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1469",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1469_ack_0,
          idata => idata,
          odata => i194x_x2_1469,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1469
    phi_stmt_1476: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1480_wire_constant & type_cast_1482_wire;
      req <= phi_stmt_1476_req_0 & phi_stmt_1476_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1476",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1476_ack_0,
          idata => idata,
          odata => k186x_x1_1476,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1476
    phi_stmt_1856: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1859_wire & type_cast_1861_wire;
      req <= phi_stmt_1856_req_0 & phi_stmt_1856_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1856",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1856_ack_0,
          idata => idata,
          odata => j240x_x0x_xph_1856,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1856
    phi_stmt_1862: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1865_wire & type_cast_1867_wire;
      req <= phi_stmt_1862_req_0 & phi_stmt_1862_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1862",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1862_ack_0,
          idata => idata,
          odata => i194x_x1x_xph_1862,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1862
    phi_stmt_1868: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1871_wire & type_cast_1874_wire_constant;
      req <= phi_stmt_1868_req_0 & phi_stmt_1868_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1868",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1868_ack_0,
          idata => idata,
          odata => k186x_x0x_xph_1868,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1868
    phi_stmt_2015: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2018_wire & type_cast_2021_wire_constant;
      req <= phi_stmt_2015_req_0 & phi_stmt_2015_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2015",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2015_ack_0,
          idata => idata,
          odata => k402x_x1_2015,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2015
    phi_stmt_2022: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2025_wire & type_cast_2027_wire;
      req <= phi_stmt_2022_req_0 & phi_stmt_2022_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2022",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2022_ack_0,
          idata => idata,
          odata => i406x_x2_2022,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2022
    phi_stmt_2028: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2031_wire & type_cast_2034_wire_constant;
      req <= phi_stmt_2028_req_0 & phi_stmt_2028_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2028",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2028_ack_0,
          idata => idata,
          odata => j456x_x1_2028,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2028
    phi_stmt_2421: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2424_wire & type_cast_2427_wire_constant;
      req <= phi_stmt_2421_req_0 & phi_stmt_2421_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2421",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2421_ack_0,
          idata => idata,
          odata => k402x_x0x_xph_2421,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2421
    phi_stmt_2428: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2431_wire & type_cast_2433_wire;
      req <= phi_stmt_2428_req_0 & phi_stmt_2428_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2428",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2428_ack_0,
          idata => idata,
          odata => i406x_x1x_xph_2428,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2428
    phi_stmt_2434: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2437_wire & type_cast_2439_wire;
      req <= phi_stmt_2434_req_0 & phi_stmt_2434_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2434",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2434_ack_0,
          idata => idata,
          odata => j456x_x0x_xph_2434,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2434
    phi_stmt_2590: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2594_wire_constant & type_cast_2596_wire;
      req <= phi_stmt_2590_req_0 & phi_stmt_2590_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2590",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2590_ack_0,
          idata => idata,
          odata => k620x_x1_2590,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2590
    phi_stmt_2597: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2600_wire & type_cast_2602_wire;
      req <= phi_stmt_2597_req_0 & phi_stmt_2597_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2597",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2597_ack_0,
          idata => idata,
          odata => i628x_x2_2597,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2597
    phi_stmt_2603: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2606_wire & type_cast_2608_wire;
      req <= phi_stmt_2603_req_0 & phi_stmt_2603_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2603",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2603_ack_0,
          idata => idata,
          odata => j678x_x1_2603,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2603
    phi_stmt_2982: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2985_wire & type_cast_2988_wire_constant;
      req <= phi_stmt_2982_req_0 & phi_stmt_2982_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2982",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2982_ack_0,
          idata => idata,
          odata => k620x_x0x_xph_2982,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2982
    phi_stmt_2989: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2992_wire & type_cast_2994_wire;
      req <= phi_stmt_2989_req_0 & phi_stmt_2989_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2989",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2989_ack_0,
          idata => idata,
          odata => i628x_x1x_xph_2989,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2989
    phi_stmt_2995: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2998_wire & type_cast_3000_wire;
      req <= phi_stmt_2995_req_0 & phi_stmt_2995_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2995",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2995_ack_0,
          idata => idata,
          odata => j678x_x0x_xph_2995,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2995
    phi_stmt_3141: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3144_wire & type_cast_3147_wire_constant;
      req <= phi_stmt_3141_req_0 & phi_stmt_3141_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3141",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3141_ack_0,
          idata => idata,
          odata => k840x_x1_3141,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3141
    phi_stmt_3148: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3151_wire & type_cast_3153_wire;
      req <= phi_stmt_3148_req_0 & phi_stmt_3148_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3148",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3148_ack_0,
          idata => idata,
          odata => i844x_x2_3148,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3148
    phi_stmt_3154: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3157_wire & type_cast_3160_wire_constant;
      req <= phi_stmt_3154_req_0 & phi_stmt_3154_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3154",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3154_ack_0,
          idata => idata,
          odata => j894x_x1_3154,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3154
    phi_stmt_3559: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3562_wire & type_cast_3565_wire_constant;
      req <= phi_stmt_3559_req_0 & phi_stmt_3559_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3559",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3559_ack_0,
          idata => idata,
          odata => k840x_x0x_xph_3559,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3559
    phi_stmt_3566: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3569_wire & type_cast_3571_wire;
      req <= phi_stmt_3566_req_0 & phi_stmt_3566_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3566",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3566_ack_0,
          idata => idata,
          odata => i844x_x1x_xph_3566,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3566
    phi_stmt_3572: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3575_wire & type_cast_3577_wire;
      req <= phi_stmt_3572_req_0 & phi_stmt_3572_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3572",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3572_ack_0,
          idata => idata,
          odata => j894x_x0x_xph_3572,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3572
    phi_stmt_3728: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3731_wire & type_cast_3734_wire_constant;
      req <= phi_stmt_3728_req_0 & phi_stmt_3728_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3728",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3728_ack_0,
          idata => idata,
          odata => k1060x_x1_3728,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3728
    phi_stmt_3735: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3738_wire & type_cast_3740_wire;
      req <= phi_stmt_3735_req_0 & phi_stmt_3735_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3735",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3735_ack_0,
          idata => idata,
          odata => i1068x_x2_3735,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3735
    phi_stmt_3741: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3744_wire & type_cast_3746_wire;
      req <= phi_stmt_3741_req_0 & phi_stmt_3741_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3741",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3741_ack_0,
          idata => idata,
          odata => j1118x_x1_3741,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3741
    phi_stmt_4132: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4135_wire & type_cast_4138_wire_constant;
      req <= phi_stmt_4132_req_0 & phi_stmt_4132_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4132",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4132_ack_0,
          idata => idata,
          odata => k1060x_x0x_xph_4132,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4132
    phi_stmt_4139: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4142_wire & type_cast_4144_wire;
      req <= phi_stmt_4139_req_0 & phi_stmt_4139_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4139",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4139_ack_0,
          idata => idata,
          odata => i1068x_x1x_xph_4139,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4139
    phi_stmt_4145: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4148_wire & type_cast_4150_wire;
      req <= phi_stmt_4145_req_0 & phi_stmt_4145_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4145",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4145_ack_0,
          idata => idata,
          odata => j1118x_x0x_xph_4145,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4145
    phi_stmt_4297: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4301_wire_constant & type_cast_4303_wire;
      req <= phi_stmt_4297_req_0 & phi_stmt_4297_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4297",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4297_ack_0,
          idata => idata,
          odata => k1282x_x1_4297,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4297
    phi_stmt_4304: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4307_wire & type_cast_4309_wire;
      req <= phi_stmt_4304_req_0 & phi_stmt_4304_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4304",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4304_ack_0,
          idata => idata,
          odata => i1286x_x2_4304,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4304
    phi_stmt_4310: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4314_wire_constant & type_cast_4316_wire;
      req <= phi_stmt_4310_req_0 & phi_stmt_4310_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4310",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4310_ack_0,
          idata => idata,
          odata => j1337x_x1_4310,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4310
    phi_stmt_4691: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4694_wire & type_cast_4697_wire_constant;
      req <= phi_stmt_4691_req_0 & phi_stmt_4691_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4691",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4691_ack_0,
          idata => idata,
          odata => k1282x_x0x_xph_4691,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4691
    phi_stmt_4698: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4701_wire & type_cast_4703_wire;
      req <= phi_stmt_4698_req_0 & phi_stmt_4698_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4698",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4698_ack_0,
          idata => idata,
          odata => i1286x_x1x_xph_4698,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4698
    phi_stmt_4704: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4707_wire & type_cast_4709_wire;
      req <= phi_stmt_4704_req_0 & phi_stmt_4704_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4704",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4704_ack_0,
          idata => idata,
          odata => j1337x_x0x_xph_4704,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4704
    phi_stmt_4866: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4870_wire_constant & type_cast_4872_wire;
      req <= phi_stmt_4866_req_0 & phi_stmt_4866_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4866",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4866_ack_0,
          idata => idata,
          odata => k1499x_x1_4866,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4866
    phi_stmt_4873: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4876_wire & type_cast_4878_wire;
      req <= phi_stmt_4873_req_0 & phi_stmt_4873_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4873",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4873_ack_0,
          idata => idata,
          odata => i1507x_x2_4873,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4873
    phi_stmt_4879: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_4882_wire & type_cast_4884_wire;
      req <= phi_stmt_4879_req_0 & phi_stmt_4879_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4879",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4879_ack_0,
          idata => idata,
          odata => j1558x_x1_4879,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4879
    phi_stmt_5246: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_5250_wire_constant & type_cast_5252_wire;
      req <= phi_stmt_5246_req_0 & phi_stmt_5246_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_5246",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_5246_ack_0,
          idata => idata,
          odata => k1499x_x0x_xph_5246,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_5246
    phi_stmt_5253: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_5256_wire & type_cast_5258_wire;
      req <= phi_stmt_5253_req_0 & phi_stmt_5253_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_5253",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_5253_ack_0,
          idata => idata,
          odata => i1507x_x1x_xph_5253,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_5253
    phi_stmt_5259: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_5262_wire & type_cast_5264_wire;
      req <= phi_stmt_5259_req_0 & phi_stmt_5259_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_5259",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_5259_ack_0,
          idata => idata,
          odata => j1558x_x0x_xph_5259,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_5259
    phi_stmt_899: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_903_wire_constant & type_cast_905_wire;
      req <= phi_stmt_899_req_0 & phi_stmt_899_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_899",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_899_ack_0,
          idata => idata,
          odata => jx_x1_899,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_899
    phi_stmt_906: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_910_wire_constant & type_cast_912_wire;
      req <= phi_stmt_906_req_0 & phi_stmt_906_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_906",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_906_ack_0,
          idata => idata,
          odata => ix_x2_906,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_906
    phi_stmt_913: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_917_wire_constant & type_cast_919_wire;
      req <= phi_stmt_913_req_0 & phi_stmt_913_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_913",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_913_ack_0,
          idata => idata,
          odata => kx_x1_913,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_913
    -- flow-through select operator MUX_1270_inst
    jx_x2_1271 <= type_cast_1268_wire_constant when (cmp160_1255(0) /=  '0') else inc_1227;
    -- flow-through select operator MUX_1819_inst
    j240x_x2_1820 <= div191_1342 when (cmp374_1805(0) /=  '0') else inc365_1783;
    -- flow-through select operator MUX_2384_inst
    j456x_x2_2385 <= type_cast_2382_wire_constant when (cmp592_2369(0) /=  '0') else inc582_2341;
    -- flow-through select operator MUX_2945_inst
    j678x_x2_2946 <= div625_2456 when (cmp812_2931(0) /=  '0') else inc803_2909;
    -- flow-through select operator MUX_3516_inst
    j894x_x2_3517 <= type_cast_3514_wire_constant when (cmp1031_3501(0) /=  '0') else inc1021_3473;
    -- flow-through select operator MUX_4089_inst
    j1118x_x2_4090 <= div1065_3594 when (cmp1253_4075(0) /=  '0') else inc1244_4053;
    -- flow-through select operator MUX_4660_inst
    j1337x_x2_4661 <= type_cast_4658_wire_constant when (cmp1472_4645(0) /=  '0') else inc1462_4617;
    -- flow-through select operator MUX_5215_inst
    j1558x_x2_5216 <= div1504_4726 when (cmp1691_5201(0) /=  '0') else inc1682_5179;
    addr_of_1073_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1073_final_reg_req_0;
      addr_of_1073_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1073_final_reg_req_1;
      addr_of_1073_final_reg_ack_1<= rack(0);
      addr_of_1073_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1073_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1072_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1156_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1156_final_reg_req_0;
      addr_of_1156_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1156_final_reg_req_1;
      addr_of_1156_final_reg_ack_1<= rack(0);
      addr_of_1156_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1156_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1155_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx131_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1181_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1181_final_reg_req_0;
      addr_of_1181_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1181_final_reg_req_1;
      addr_of_1181_final_reg_ack_1<= rack(0);
      addr_of_1181_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1181_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1180_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx136_1182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1629_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1629_final_reg_req_0;
      addr_of_1629_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1629_final_reg_req_1;
      addr_of_1629_final_reg_ack_1<= rack(0);
      addr_of_1629_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1629_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1628_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx299_1630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1712_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1712_final_reg_req_0;
      addr_of_1712_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1712_final_reg_req_1;
      addr_of_1712_final_reg_ack_1<= rack(0);
      addr_of_1712_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1712_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1711_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx342_1713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1737_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1737_final_reg_req_0;
      addr_of_1737_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1737_final_reg_req_1;
      addr_of_1737_final_reg_ack_1<= rack(0);
      addr_of_1737_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1737_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1736_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx347_1738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2187_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2187_final_reg_req_0;
      addr_of_2187_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2187_final_reg_req_1;
      addr_of_2187_final_reg_ack_1<= rack(0);
      addr_of_2187_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2187_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2186_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx516_2188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2270_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2270_final_reg_req_0;
      addr_of_2270_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2270_final_reg_req_1;
      addr_of_2270_final_reg_ack_1<= rack(0);
      addr_of_2270_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2270_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2269_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx559_2271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2295_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2295_final_reg_req_0;
      addr_of_2295_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2295_final_reg_req_1;
      addr_of_2295_final_reg_ack_1<= rack(0);
      addr_of_2295_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2295_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2294_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx564_2296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2755_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2755_final_reg_req_0;
      addr_of_2755_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2755_final_reg_req_1;
      addr_of_2755_final_reg_ack_1<= rack(0);
      addr_of_2755_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2755_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2754_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx737_2756,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2838_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2838_final_reg_req_0;
      addr_of_2838_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2838_final_reg_req_1;
      addr_of_2838_final_reg_ack_1<= rack(0);
      addr_of_2838_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2838_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2837_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx780_2839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2863_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2863_final_reg_req_0;
      addr_of_2863_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2863_final_reg_req_1;
      addr_of_2863_final_reg_ack_1<= rack(0);
      addr_of_2863_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2863_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2862_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx785_2864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3319_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3319_final_reg_req_0;
      addr_of_3319_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3319_final_reg_req_1;
      addr_of_3319_final_reg_ack_1<= rack(0);
      addr_of_3319_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3319_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3318_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx955_3320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3402_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3402_final_reg_req_0;
      addr_of_3402_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3402_final_reg_req_1;
      addr_of_3402_final_reg_ack_1<= rack(0);
      addr_of_3402_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3402_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3401_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx998_3403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3427_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3427_final_reg_req_0;
      addr_of_3427_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3427_final_reg_req_1;
      addr_of_3427_final_reg_ack_1<= rack(0);
      addr_of_3427_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3427_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3426_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1003_3428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3899_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3899_final_reg_req_0;
      addr_of_3899_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3899_final_reg_req_1;
      addr_of_3899_final_reg_ack_1<= rack(0);
      addr_of_3899_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3899_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3898_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1178_3900,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3982_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3982_final_reg_req_0;
      addr_of_3982_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3982_final_reg_req_1;
      addr_of_3982_final_reg_ack_1<= rack(0);
      addr_of_3982_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3982_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3981_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1221_3983,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4007_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4007_final_reg_req_0;
      addr_of_4007_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4007_final_reg_req_1;
      addr_of_4007_final_reg_ack_1<= rack(0);
      addr_of_4007_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4007_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4006_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1226_4008,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4463_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4463_final_reg_req_0;
      addr_of_4463_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4463_final_reg_req_1;
      addr_of_4463_final_reg_ack_1<= rack(0);
      addr_of_4463_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4463_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4462_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1396_4464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4546_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4546_final_reg_req_0;
      addr_of_4546_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4546_final_reg_req_1;
      addr_of_4546_final_reg_ack_1<= rack(0);
      addr_of_4546_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4546_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4545_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1439_4547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_4571_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_4571_final_reg_req_0;
      addr_of_4571_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_4571_final_reg_req_1;
      addr_of_4571_final_reg_ack_1<= rack(0);
      addr_of_4571_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_4571_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_4570_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1444_4572,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_5025_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_5025_final_reg_req_0;
      addr_of_5025_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_5025_final_reg_req_1;
      addr_of_5025_final_reg_ack_1<= rack(0);
      addr_of_5025_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_5025_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_5024_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1616_5026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_5108_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_5108_final_reg_req_0;
      addr_of_5108_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_5108_final_reg_req_1;
      addr_of_5108_final_reg_ack_1<= rack(0);
      addr_of_5108_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_5108_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_5107_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1659_5109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_5133_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_5133_final_reg_req_0;
      addr_of_5133_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_5133_final_reg_req_1;
      addr_of_5133_final_reg_ack_1<= rack(0);
      addr_of_5133_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_5133_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_5132_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1664_5134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1011_inst
    process(conv60_976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv60_976(31 downto 0);
      type_cast_1011_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1013_inst
    process(add73_1008) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add73_1008(31 downto 0);
      type_cast_1013_wire <= tmp_var; -- 
    end process;
    type_cast_1026_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1026_inst_req_0;
      type_cast_1026_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1026_inst_req_1;
      type_cast_1026_inst_ack_1<= rack(0);
      type_cast_1026_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1026_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1025_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_1027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1031_inst_req_0;
      type_cast_1031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1031_inst_req_1;
      type_cast_1031_inst_ack_1<= rack(0);
      type_cast_1031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1030_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1055_inst
    process(add90_1052) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add90_1052(31 downto 0);
      type_cast_1055_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1060_inst
    process(ASHR_i32_i32_1059_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1059_wire(31 downto 0);
      shr_1061 <= tmp_var; -- 
    end process;
    type_cast_1066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1066_inst_req_0;
      type_cast_1066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1066_inst_req_1;
      type_cast_1066_inst_ack_1<= rack(0);
      type_cast_1066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1065_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1067,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1085_inst_req_0;
      type_cast_1085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1085_inst_req_1;
      type_cast_1085_inst_ack_1<= rack(0);
      type_cast_1085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1084_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1086,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1139_inst
    process(add111_1116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add111_1116(31 downto 0);
      type_cast_1139_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1144_inst
    process(ASHR_i32_i32_1143_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1143_wire(31 downto 0);
      shr129_1145 <= tmp_var; -- 
    end process;
    type_cast_1149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1149_inst_req_0;
      type_cast_1149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1149_inst_req_1;
      type_cast_1149_inst_ack_1<= rack(0);
      type_cast_1149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1148_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom130_1150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1164_inst
    process(add127_1136) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add127_1136(31 downto 0);
      type_cast_1164_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1169_inst
    process(ASHR_i32_i32_1168_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1168_wire(31 downto 0);
      shr134_1170 <= tmp_var; -- 
    end process;
    type_cast_1174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1174_inst_req_0;
      type_cast_1174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1174_inst_req_1;
      type_cast_1174_inst_ack_1<= rack(0);
      type_cast_1174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1173_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom135_1175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1192_inst_req_0;
      type_cast_1192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1192_inst_req_1;
      type_cast_1192_inst_ack_1<= rack(0);
      type_cast_1192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1191_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv139_1193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1202_inst
    process(add140_1199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add140_1199(31 downto 0);
      type_cast_1202_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1204_inst
    process(conv31_811) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv31_811(31 downto 0);
      type_cast_1204_wire <= tmp_var; -- 
    end process;
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack(0);
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1230_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp154_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1258_inst_req_0;
      type_cast_1258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1258_inst_req_1;
      type_cast_1258_inst_ack_1<= rack(0);
      type_cast_1258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp160_1255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc165_1259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1275_inst_req_0;
      type_cast_1275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1275_inst_req_1;
      type_cast_1275_inst_ack_1<= rack(0);
      type_cast_1275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1274_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv168_1276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1282_inst_req_0;
      type_cast_1282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1282_inst_req_1;
      type_cast_1282_inst_ack_1<= rack(0);
      type_cast_1282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp169_1279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1310_inst_req_0;
      type_cast_1310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1310_inst_req_1;
      type_cast_1310_inst_ack_1<= rack(0);
      type_cast_1310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1310_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1312_inst_req_0;
      type_cast_1312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1312_inst_req_1;
      type_cast_1312_inst_ack_1<= rack(0);
      type_cast_1312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_899,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1312_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1316_inst_req_0;
      type_cast_1316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1316_inst_req_1;
      type_cast_1316_inst_ack_1<= rack(0);
      type_cast_1316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1316_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1318_inst_req_0;
      type_cast_1318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1318_inst_req_1;
      type_cast_1318_inst_ack_1<= rack(0);
      type_cast_1318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc165x_xix_x2_1264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1318_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1325_inst_req_0;
      type_cast_1325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1325_inst_req_1;
      type_cast_1325_inst_ack_1<= rack(0);
      type_cast_1325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add148_1219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1325_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1335_inst_req_0;
      type_cast_1335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1335_inst_req_1;
      type_cast_1335_inst_ack_1<= rack(0);
      type_cast_1335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp189_1332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv190_1336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1375_inst_req_0;
      type_cast_1375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1375_inst_req_1;
      type_cast_1375_inst_ack_1<= rack(0);
      type_cast_1375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp201_1348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv226_1376,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1379_inst_req_0;
      type_cast_1379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1379_inst_req_1;
      type_cast_1379_inst_ack_1<= rack(0);
      type_cast_1379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1379_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp189_1332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv228_1380,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1389_inst
    process(sext1766_1386) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1766_1386(31 downto 0);
      type_cast_1389_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1394_inst
    process(ASHR_i32_i32_1393_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1393_wire(31 downto 0);
      conv234_1395 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1404_inst
    process(sext1718_1401) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1718_1401(31 downto 0);
      type_cast_1404_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1409_inst
    process(ASHR_i32_i32_1408_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1408_wire(31 downto 0);
      conv236_1410 <= tmp_var; -- 
    end process;
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp197_1345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv248_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1428_inst
    process(sext1767_1425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1767_1425(31 downto 0);
      type_cast_1428_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1433_inst
    process(ASHR_i32_i32_1432_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1432_wire(31 downto 0);
      conv291_1434 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1454_inst
    process(sext1719_1451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1719_1451(31 downto 0);
      type_cast_1454_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1459_inst
    process(ASHR_i32_i32_1458_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1458_wire(31 downto 0);
      conv315_1460 <= tmp_var; -- 
    end process;
    type_cast_1466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1466_inst_req_0;
      type_cast_1466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1466_inst_req_1;
      type_cast_1466_inst_ack_1<= rack(0);
      type_cast_1466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div191_1342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1466_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1468_inst_req_0;
      type_cast_1468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1468_inst_req_1;
      type_cast_1468_inst_ack_1<= rack(0);
      type_cast_1468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j240x_x0x_xph_1856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1468_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1475_inst_req_0;
      type_cast_1475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1475_inst_req_1;
      type_cast_1475_inst_ack_1<= rack(0);
      type_cast_1475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i194x_x1x_xph_1862,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1475_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1482_inst_req_0;
      type_cast_1482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1482_inst_req_1;
      type_cast_1482_inst_ack_1<= rack(0);
      type_cast_1482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k186x_x0x_xph_1868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1482_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1487_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1487_inst_req_0;
      type_cast_1487_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1487_inst_req_1;
      type_cast_1487_inst_ack_1<= rack(0);
      type_cast_1487_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1487_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1486_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv246_1488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1491_inst
    process(conv246_1488) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv246_1488(31 downto 0);
      type_cast_1491_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1493_inst
    process(conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv248_1419(31 downto 0);
      type_cast_1493_wire <= tmp_var; -- 
    end process;
    type_cast_1508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1508_inst_req_0;
      type_cast_1508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1508_inst_req_1;
      type_cast_1508_inst_ack_1<= rack(0);
      type_cast_1508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp254_1505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1523_inst
    process(conv246_1488) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv246_1488(31 downto 0);
      type_cast_1523_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1525_inst
    process(add259_1520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add259_1520(31 downto 0);
      type_cast_1525_wire <= tmp_var; -- 
    end process;
    type_cast_1538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1538_inst_req_0;
      type_cast_1538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1538_inst_req_1;
      type_cast_1538_inst_ack_1<= rack(0);
      type_cast_1538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1537_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv264_1539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1542_inst
    process(conv264_1539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv264_1539(31 downto 0);
      type_cast_1542_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1544_inst
    process(conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv248_1419(31 downto 0);
      type_cast_1544_wire <= tmp_var; -- 
    end process;
    type_cast_1559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1559_inst_req_0;
      type_cast_1559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1559_inst_req_1;
      type_cast_1559_inst_ack_1<= rack(0);
      type_cast_1559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp272_1556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv273_1560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1568_inst
    process(conv264_1539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv264_1539(31 downto 0);
      type_cast_1568_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1570_inst
    process(add276_1565) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add276_1565(31 downto 0);
      type_cast_1570_wire <= tmp_var; -- 
    end process;
    type_cast_1583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1583_inst_req_0;
      type_cast_1583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1583_inst_req_1;
      type_cast_1583_inst_ack_1<= rack(0);
      type_cast_1583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1582_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv283_1584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1588_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1588_inst_req_0;
      type_cast_1588_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1588_inst_req_1;
      type_cast_1588_inst_ack_1<= rack(0);
      type_cast_1588_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1588_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1587_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv287_1589,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1612_inst
    process(add295_1609) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add295_1609(31 downto 0);
      type_cast_1612_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1617_inst
    process(ASHR_i32_i32_1616_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1616_wire(31 downto 0);
      shr297_1618 <= tmp_var; -- 
    end process;
    type_cast_1622_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1622_inst_req_0;
      type_cast_1622_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1622_inst_req_1;
      type_cast_1622_inst_ack_1<= rack(0);
      type_cast_1622_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1622_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1621_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom298_1623,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1641_inst_req_0;
      type_cast_1641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1641_inst_req_1;
      type_cast_1641_inst_ack_1<= rack(0);
      type_cast_1641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1641_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1640_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_1642,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1695_inst
    process(add322_1672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add322_1672(31 downto 0);
      type_cast_1695_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1700_inst
    process(ASHR_i32_i32_1699_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1699_wire(31 downto 0);
      shr340_1701 <= tmp_var; -- 
    end process;
    type_cast_1705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1705_inst_req_0;
      type_cast_1705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1705_inst_req_1;
      type_cast_1705_inst_ack_1<= rack(0);
      type_cast_1705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1704_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom341_1706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1720_inst
    process(add338_1692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add338_1692(31 downto 0);
      type_cast_1720_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1725_inst
    process(ASHR_i32_i32_1724_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1724_wire(31 downto 0);
      shr345_1726 <= tmp_var; -- 
    end process;
    type_cast_1730_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1730_inst_req_0;
      type_cast_1730_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1730_inst_req_1;
      type_cast_1730_inst_ack_1<= rack(0);
      type_cast_1730_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1730_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1729_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom346_1731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1748_inst_req_0;
      type_cast_1748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1748_inst_req_1;
      type_cast_1748_inst_ack_1<= rack(0);
      type_cast_1748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1747_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv352_1749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1758_inst
    process(add353_1755) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add353_1755(31 downto 0);
      type_cast_1758_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1760_inst
    process(conv226_1376) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv226_1376(31 downto 0);
      type_cast_1760_wire <= tmp_var; -- 
    end process;
    type_cast_1787_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1787_inst_req_0;
      type_cast_1787_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1787_inst_req_1;
      type_cast_1787_inst_ack_1<= rack(0);
      type_cast_1787_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1787_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1786_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1794_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1794_inst_req_0;
      type_cast_1794_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1794_inst_req_1;
      type_cast_1794_inst_ack_1<= rack(0);
      type_cast_1794_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1794_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp368_1791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv369_1795,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1808_inst_req_0;
      type_cast_1808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1808_inst_req_1;
      type_cast_1808_inst_ack_1<= rack(0);
      type_cast_1808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp374_1805,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc379_1809,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1824_inst_req_0;
      type_cast_1824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1824_inst_req_1;
      type_cast_1824_inst_ack_1<= rack(0);
      type_cast_1824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1823_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv382_1825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1831_inst_req_0;
      type_cast_1831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1831_inst_req_1;
      type_cast_1831_inst_ack_1<= rack(0);
      type_cast_1831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp383_1828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv384_1832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1859_inst_req_0;
      type_cast_1859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1859_inst_req_1;
      type_cast_1859_inst_ack_1<= rack(0);
      type_cast_1859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j240x_x1_1463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1859_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1861_inst_req_0;
      type_cast_1861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1861_inst_req_1;
      type_cast_1861_inst_ack_1<= rack(0);
      type_cast_1861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j240x_x2_1820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1861_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1865_inst_req_0;
      type_cast_1865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1865_inst_req_1;
      type_cast_1865_inst_ack_1<= rack(0);
      type_cast_1865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i194x_x2_1469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1865_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1867_inst_req_0;
      type_cast_1867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1867_inst_req_1;
      type_cast_1867_inst_ack_1<= rack(0);
      type_cast_1867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1867_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc379x_xi194x_x2_1814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1867_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1871_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1871_inst_req_0;
      type_cast_1871_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1871_inst_req_1;
      type_cast_1871_inst_ack_1<= rack(0);
      type_cast_1871_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1871_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add361_1775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1871_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1884_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1884_inst_req_0;
      type_cast_1884_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1884_inst_req_1;
      type_cast_1884_inst_ack_1<= rack(0);
      type_cast_1884_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1884_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp407_1881,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv408_1885,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1927_inst_req_0;
      type_cast_1927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1927_inst_req_1;
      type_cast_1927_inst_ack_1<= rack(0);
      type_cast_1927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp417_1897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv442_1928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1931_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1931_inst_req_0;
      type_cast_1931_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1931_inst_req_1;
      type_cast_1931_inst_ack_1<= rack(0);
      type_cast_1931_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1931_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp421_1900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv444_1932,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1941_inst
    process(sext1768_1938) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1768_1938(31 downto 0);
      type_cast_1941_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1946_inst
    process(ASHR_i32_i32_1945_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1945_wire(31 downto 0);
      conv450_1947 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1956_inst
    process(sext1720_1953) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1720_1953(31 downto 0);
      type_cast_1956_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1961_inst
    process(ASHR_i32_i32_1960_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1960_wire(31 downto 0);
      conv452_1962 <= tmp_var; -- 
    end process;
    type_cast_1970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1970_inst_req_0;
      type_cast_1970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1970_inst_req_1;
      type_cast_1970_inst_ack_1<= rack(0);
      type_cast_1970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp413_1894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv464_1971,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1980_inst
    process(sext1769_1977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1769_1977(31 downto 0);
      type_cast_1980_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1985_inst
    process(ASHR_i32_i32_1984_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1984_wire(31 downto 0);
      conv508_1986 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2006_inst
    process(sext1721_2003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1721_2003(31 downto 0);
      type_cast_2006_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2011_inst
    process(ASHR_i32_i32_2010_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2010_wire(31 downto 0);
      conv532_2012 <= tmp_var; -- 
    end process;
    type_cast_2018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2018_inst_req_0;
      type_cast_2018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2018_inst_req_1;
      type_cast_2018_inst_ack_1<= rack(0);
      type_cast_2018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k402x_x0x_xph_2421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2018_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2025_inst_req_0;
      type_cast_2025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2025_inst_req_1;
      type_cast_2025_inst_ack_1<= rack(0);
      type_cast_2025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div409_1891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2025_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2027_inst_req_0;
      type_cast_2027_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2027_inst_req_1;
      type_cast_2027_inst_ack_1<= rack(0);
      type_cast_2027_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2027_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i406x_x1x_xph_2428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2027_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2031_inst_req_0;
      type_cast_2031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2031_inst_req_1;
      type_cast_2031_inst_ack_1<= rack(0);
      type_cast_2031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j456x_x0x_xph_2434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2031_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2039_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2039_inst_req_0;
      type_cast_2039_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2039_inst_req_1;
      type_cast_2039_inst_ack_1<= rack(0);
      type_cast_2039_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2039_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2038_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv462_2040,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2043_inst
    process(conv462_2040) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv462_2040(31 downto 0);
      type_cast_2043_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2045_inst
    process(conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv464_1971(31 downto 0);
      type_cast_2045_wire <= tmp_var; -- 
    end process;
    type_cast_2060_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2060_inst_req_0;
      type_cast_2060_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2060_inst_req_1;
      type_cast_2060_inst_ack_1<= rack(0);
      type_cast_2060_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2060_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp470_2057,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv471_2061,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2075_inst
    process(conv462_2040) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv462_2040(31 downto 0);
      type_cast_2075_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2077_inst
    process(add475_2072) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add475_2072(31 downto 0);
      type_cast_2077_wire <= tmp_var; -- 
    end process;
    type_cast_2090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2090_inst_req_0;
      type_cast_2090_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2090_inst_req_1;
      type_cast_2090_inst_ack_1<= rack(0);
      type_cast_2090_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2090_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2089_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv480_2091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2094_inst
    process(conv480_2091) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv480_2091(31 downto 0);
      type_cast_2094_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2096_inst
    process(conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv464_1971(31 downto 0);
      type_cast_2096_wire <= tmp_var; -- 
    end process;
    type_cast_2111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2111_inst_req_0;
      type_cast_2111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2111_inst_req_1;
      type_cast_2111_inst_ack_1<= rack(0);
      type_cast_2111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp488_2108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv489_2112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2126_inst
    process(conv480_2091) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv480_2091(31 downto 0);
      type_cast_2126_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2128_inst
    process(add493_2123) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add493_2123(31 downto 0);
      type_cast_2128_wire <= tmp_var; -- 
    end process;
    type_cast_2141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2141_inst_req_0;
      type_cast_2141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2141_inst_req_1;
      type_cast_2141_inst_ack_1<= rack(0);
      type_cast_2141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2140_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv500_2142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2146_inst_req_0;
      type_cast_2146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2146_inst_req_1;
      type_cast_2146_inst_ack_1<= rack(0);
      type_cast_2146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2145_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv504_2147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2170_inst
    process(add512_2167) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add512_2167(31 downto 0);
      type_cast_2170_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2175_inst
    process(ASHR_i32_i32_2174_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2174_wire(31 downto 0);
      shr514_2176 <= tmp_var; -- 
    end process;
    type_cast_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2180_inst_req_0;
      type_cast_2180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2180_inst_req_1;
      type_cast_2180_inst_ack_1<= rack(0);
      type_cast_2180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2179_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom515_2181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2198_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv521_2200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2253_inst
    process(add539_2230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add539_2230(31 downto 0);
      type_cast_2253_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2258_inst
    process(ASHR_i32_i32_2257_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2257_wire(31 downto 0);
      shr557_2259 <= tmp_var; -- 
    end process;
    type_cast_2263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2263_inst_req_0;
      type_cast_2263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2263_inst_req_1;
      type_cast_2263_inst_ack_1<= rack(0);
      type_cast_2263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2262_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom558_2264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2278_inst
    process(add555_2250) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add555_2250(31 downto 0);
      type_cast_2278_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2283_inst
    process(ASHR_i32_i32_2282_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2282_wire(31 downto 0);
      shr562_2284 <= tmp_var; -- 
    end process;
    type_cast_2288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2288_inst_req_0;
      type_cast_2288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2288_inst_req_1;
      type_cast_2288_inst_ack_1<= rack(0);
      type_cast_2288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2287_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom563_2289,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2306_inst_req_0;
      type_cast_2306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2306_inst_req_1;
      type_cast_2306_inst_ack_1<= rack(0);
      type_cast_2306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2305_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv569_2307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2316_inst
    process(add570_2313) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add570_2313(31 downto 0);
      type_cast_2316_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2318_inst
    process(conv442_1928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv442_1928(31 downto 0);
      type_cast_2318_wire <= tmp_var; -- 
    end process;
    type_cast_2345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2345_inst_req_0;
      type_cast_2345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2345_inst_req_1;
      type_cast_2345_inst_ack_1<= rack(0);
      type_cast_2345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2344_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv584_2346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2352_inst_req_0;
      type_cast_2352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2352_inst_req_1;
      type_cast_2352_inst_ack_1<= rack(0);
      type_cast_2352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp585_2349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv586_2353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2372_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2372_inst_req_0;
      type_cast_2372_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2372_inst_req_1;
      type_cast_2372_inst_ack_1<= rack(0);
      type_cast_2372_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2372_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp592_2369,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc597_2373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2389_inst_req_0;
      type_cast_2389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2389_inst_req_1;
      type_cast_2389_inst_ack_1<= rack(0);
      type_cast_2389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2388_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv600_2390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2396_inst_req_0;
      type_cast_2396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2396_inst_req_1;
      type_cast_2396_inst_ack_1<= rack(0);
      type_cast_2396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp601_2393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv602_2397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2424_inst_req_0;
      type_cast_2424_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2424_inst_req_1;
      type_cast_2424_inst_ack_1<= rack(0);
      type_cast_2424_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2424_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add578_2333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2424_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2431_inst_req_0;
      type_cast_2431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2431_inst_req_1;
      type_cast_2431_inst_ack_1<= rack(0);
      type_cast_2431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i406x_x2_2022,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2431_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2433_inst_req_0;
      type_cast_2433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2433_inst_req_1;
      type_cast_2433_inst_ack_1<= rack(0);
      type_cast_2433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc597x_xi406x_x2_2378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2433_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2437_inst_req_0;
      type_cast_2437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2437_inst_req_1;
      type_cast_2437_inst_ack_1<= rack(0);
      type_cast_2437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j456x_x1_2028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2437_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2439_inst_req_0;
      type_cast_2439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2439_inst_req_1;
      type_cast_2439_inst_ack_1<= rack(0);
      type_cast_2439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j456x_x2_2385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2439_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2449_inst_req_0;
      type_cast_2449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2449_inst_req_1;
      type_cast_2449_inst_ack_1<= rack(0);
      type_cast_2449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp623_2446,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv624_2450,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2462_inst_req_0;
      type_cast_2462_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2462_inst_req_1;
      type_cast_2462_inst_ack_1<= rack(0);
      type_cast_2462_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2462_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp629_2459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv630_2463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2502_inst_req_0;
      type_cast_2502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2502_inst_req_1;
      type_cast_2502_inst_ack_1<= rack(0);
      type_cast_2502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp639_2475,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv664_2503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2506_inst_req_0;
      type_cast_2506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2506_inst_req_1;
      type_cast_2506_inst_ack_1<= rack(0);
      type_cast_2506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp623_2446,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv666_2507,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2516_inst
    process(sext1770_2513) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1770_2513(31 downto 0);
      type_cast_2516_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2521_inst
    process(ASHR_i32_i32_2520_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2520_wire(31 downto 0);
      conv672_2522 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2531_inst
    process(sext1722_2528) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1722_2528(31 downto 0);
      type_cast_2531_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2536_inst
    process(ASHR_i32_i32_2535_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2535_wire(31 downto 0);
      conv674_2537 <= tmp_var; -- 
    end process;
    type_cast_2545_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2545_inst_req_0;
      type_cast_2545_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2545_inst_req_1;
      type_cast_2545_inst_ack_1<= rack(0);
      type_cast_2545_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2545_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp635_2472,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv686_2546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2555_inst
    process(sext1771_2552) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1771_2552(31 downto 0);
      type_cast_2555_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2560_inst
    process(ASHR_i32_i32_2559_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2559_wire(31 downto 0);
      conv729_2561 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2581_inst
    process(sext1723_2578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1723_2578(31 downto 0);
      type_cast_2581_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2586_inst
    process(ASHR_i32_i32_2585_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2585_wire(31 downto 0);
      conv753_2587 <= tmp_var; -- 
    end process;
    type_cast_2596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2596_inst_req_0;
      type_cast_2596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2596_inst_req_1;
      type_cast_2596_inst_ack_1<= rack(0);
      type_cast_2596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k620x_x0x_xph_2982,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2596_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2600_inst_req_0;
      type_cast_2600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2600_inst_req_1;
      type_cast_2600_inst_ack_1<= rack(0);
      type_cast_2600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div631_2469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2600_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2602_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2602_inst_req_0;
      type_cast_2602_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2602_inst_req_1;
      type_cast_2602_inst_ack_1<= rack(0);
      type_cast_2602_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2602_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i628x_x1x_xph_2989,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2602_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2606_inst_req_0;
      type_cast_2606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2606_inst_req_1;
      type_cast_2606_inst_ack_1<= rack(0);
      type_cast_2606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div625_2456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2606_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2608_inst_req_0;
      type_cast_2608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2608_inst_req_1;
      type_cast_2608_inst_ack_1<= rack(0);
      type_cast_2608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j678x_x0x_xph_2995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2608_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2613_inst_req_0;
      type_cast_2613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2613_inst_req_1;
      type_cast_2613_inst_ack_1<= rack(0);
      type_cast_2613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2612_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv684_2614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2617_inst
    process(conv684_2614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv684_2614(31 downto 0);
      type_cast_2617_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2619_inst
    process(conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv686_2546(31 downto 0);
      type_cast_2619_wire <= tmp_var; -- 
    end process;
    type_cast_2634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2634_inst_req_0;
      type_cast_2634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2634_inst_req_1;
      type_cast_2634_inst_ack_1<= rack(0);
      type_cast_2634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp692_2631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv693_2635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2649_inst
    process(conv684_2614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv684_2614(31 downto 0);
      type_cast_2649_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2651_inst
    process(add697_2646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add697_2646(31 downto 0);
      type_cast_2651_wire <= tmp_var; -- 
    end process;
    type_cast_2664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2664_inst_req_0;
      type_cast_2664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2664_inst_req_1;
      type_cast_2664_inst_ack_1<= rack(0);
      type_cast_2664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2663_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv702_2665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2668_inst
    process(conv702_2665) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv702_2665(31 downto 0);
      type_cast_2668_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2670_inst
    process(conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv686_2546(31 downto 0);
      type_cast_2670_wire <= tmp_var; -- 
    end process;
    type_cast_2685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2685_inst_req_0;
      type_cast_2685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2685_inst_req_1;
      type_cast_2685_inst_ack_1<= rack(0);
      type_cast_2685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp710_2682,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv711_2686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2694_inst
    process(conv702_2665) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv702_2665(31 downto 0);
      type_cast_2694_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2696_inst
    process(add714_2691) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add714_2691(31 downto 0);
      type_cast_2696_wire <= tmp_var; -- 
    end process;
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2708_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv721_2710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2714_inst_req_0;
      type_cast_2714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2714_inst_req_1;
      type_cast_2714_inst_ack_1<= rack(0);
      type_cast_2714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2713_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv725_2715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2738_inst
    process(add733_2735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add733_2735(31 downto 0);
      type_cast_2738_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2743_inst
    process(ASHR_i32_i32_2742_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2742_wire(31 downto 0);
      shr735_2744 <= tmp_var; -- 
    end process;
    type_cast_2748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2748_inst_req_0;
      type_cast_2748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2748_inst_req_1;
      type_cast_2748_inst_ack_1<= rack(0);
      type_cast_2748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2747_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom736_2749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2767_inst_req_0;
      type_cast_2767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2767_inst_req_1;
      type_cast_2767_inst_ack_1<= rack(0);
      type_cast_2767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2766_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv742_2768,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2821_inst
    process(add760_2798) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add760_2798(31 downto 0);
      type_cast_2821_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2826_inst
    process(ASHR_i32_i32_2825_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2825_wire(31 downto 0);
      shr778_2827 <= tmp_var; -- 
    end process;
    type_cast_2831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2831_inst_req_0;
      type_cast_2831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2831_inst_req_1;
      type_cast_2831_inst_ack_1<= rack(0);
      type_cast_2831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2830_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom779_2832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2846_inst
    process(add776_2818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add776_2818(31 downto 0);
      type_cast_2846_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2851_inst
    process(ASHR_i32_i32_2850_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2850_wire(31 downto 0);
      shr783_2852 <= tmp_var; -- 
    end process;
    type_cast_2856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2856_inst_req_0;
      type_cast_2856_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2856_inst_req_1;
      type_cast_2856_inst_ack_1<= rack(0);
      type_cast_2856_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2856_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2855_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom784_2857,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2874_inst_req_0;
      type_cast_2874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2874_inst_req_1;
      type_cast_2874_inst_ack_1<= rack(0);
      type_cast_2874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2873_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv790_2875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2884_inst
    process(add791_2881) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add791_2881(31 downto 0);
      type_cast_2884_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2886_inst
    process(conv664_2503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv664_2503(31 downto 0);
      type_cast_2886_wire <= tmp_var; -- 
    end process;
    type_cast_2913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2913_inst_req_0;
      type_cast_2913_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2913_inst_req_1;
      type_cast_2913_inst_ack_1<= rack(0);
      type_cast_2913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2913_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2912_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv805_2914,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2920_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2920_inst_req_0;
      type_cast_2920_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2920_inst_req_1;
      type_cast_2920_inst_ack_1<= rack(0);
      type_cast_2920_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2920_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp806_2917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv807_2921,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2934_inst_req_0;
      type_cast_2934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2934_inst_req_1;
      type_cast_2934_inst_ack_1<= rack(0);
      type_cast_2934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp812_2931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc817_2935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2950_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2950_inst_req_0;
      type_cast_2950_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2950_inst_req_1;
      type_cast_2950_inst_ack_1<= rack(0);
      type_cast_2950_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2950_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2949_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv820_2951,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2957_inst_req_0;
      type_cast_2957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2957_inst_req_1;
      type_cast_2957_inst_ack_1<= rack(0);
      type_cast_2957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp821_2954,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv822_2958,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2985_inst_req_0;
      type_cast_2985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2985_inst_req_1;
      type_cast_2985_inst_ack_1<= rack(0);
      type_cast_2985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add799_2901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2985_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2992_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2992_inst_req_0;
      type_cast_2992_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2992_inst_req_1;
      type_cast_2992_inst_ack_1<= rack(0);
      type_cast_2992_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2992_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i628x_x2_2597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2992_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2994_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2994_inst_req_0;
      type_cast_2994_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2994_inst_req_1;
      type_cast_2994_inst_ack_1<= rack(0);
      type_cast_2994_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2994_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc817x_xi628x_x2_2940,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2994_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2998_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2998_inst_req_0;
      type_cast_2998_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2998_inst_req_1;
      type_cast_2998_inst_ack_1<= rack(0);
      type_cast_2998_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2998_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j678x_x1_2603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2998_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3000_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3000_inst_req_0;
      type_cast_3000_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3000_inst_req_1;
      type_cast_3000_inst_ack_1<= rack(0);
      type_cast_3000_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3000_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j678x_x2_2946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3000_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3010_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3010_inst_req_0;
      type_cast_3010_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3010_inst_req_1;
      type_cast_3010_inst_ack_1<= rack(0);
      type_cast_3010_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3010_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp845_3007,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv846_3011,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3053_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3053_inst_req_0;
      type_cast_3053_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3053_inst_req_1;
      type_cast_3053_inst_ack_1<= rack(0);
      type_cast_3053_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3053_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp855_3023,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv880_3054,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3057_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3057_inst_req_0;
      type_cast_3057_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3057_inst_req_1;
      type_cast_3057_inst_ack_1<= rack(0);
      type_cast_3057_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3057_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp859_3026,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv882_3058,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3067_inst
    process(sext1772_3064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1772_3064(31 downto 0);
      type_cast_3067_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3072_inst
    process(ASHR_i32_i32_3071_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3071_wire(31 downto 0);
      conv888_3073 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3082_inst
    process(sext1724_3079) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1724_3079(31 downto 0);
      type_cast_3082_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3087_inst
    process(ASHR_i32_i32_3086_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3086_wire(31 downto 0);
      conv890_3088 <= tmp_var; -- 
    end process;
    type_cast_3096_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3096_inst_req_0;
      type_cast_3096_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3096_inst_req_1;
      type_cast_3096_inst_ack_1<= rack(0);
      type_cast_3096_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3096_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp851_3020,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv902_3097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3106_inst
    process(sext1773_3103) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1773_3103(31 downto 0);
      type_cast_3106_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3111_inst
    process(ASHR_i32_i32_3110_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3110_wire(31 downto 0);
      conv947_3112 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3132_inst
    process(sext1725_3129) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1725_3129(31 downto 0);
      type_cast_3132_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3137_inst
    process(ASHR_i32_i32_3136_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3136_wire(31 downto 0);
      conv971_3138 <= tmp_var; -- 
    end process;
    type_cast_3144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3144_inst_req_0;
      type_cast_3144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3144_inst_req_1;
      type_cast_3144_inst_ack_1<= rack(0);
      type_cast_3144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k840x_x0x_xph_3559,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3144_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3151_inst_req_0;
      type_cast_3151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3151_inst_req_1;
      type_cast_3151_inst_ack_1<= rack(0);
      type_cast_3151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div847_3017,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3151_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3153_inst_req_0;
      type_cast_3153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3153_inst_req_1;
      type_cast_3153_inst_ack_1<= rack(0);
      type_cast_3153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i844x_x1x_xph_3566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3157_inst_req_0;
      type_cast_3157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3157_inst_req_1;
      type_cast_3157_inst_ack_1<= rack(0);
      type_cast_3157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j894x_x0x_xph_3572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3157_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3165_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3165_inst_req_0;
      type_cast_3165_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3165_inst_req_1;
      type_cast_3165_inst_ack_1<= rack(0);
      type_cast_3165_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3165_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3164_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv900_3166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3169_inst
    process(conv900_3166) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv900_3166(31 downto 0);
      type_cast_3169_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3171_inst
    process(conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv902_3097(31 downto 0);
      type_cast_3171_wire <= tmp_var; -- 
    end process;
    type_cast_3186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3186_inst_req_0;
      type_cast_3186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3186_inst_req_1;
      type_cast_3186_inst_ack_1<= rack(0);
      type_cast_3186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp908_3183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv909_3187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3207_inst
    process(conv900_3166) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv900_3166(31 downto 0);
      type_cast_3207_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3209_inst
    process(add914_3204) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add914_3204(31 downto 0);
      type_cast_3209_wire <= tmp_var; -- 
    end process;
    type_cast_3222_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3222_inst_req_0;
      type_cast_3222_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3222_inst_req_1;
      type_cast_3222_inst_ack_1<= rack(0);
      type_cast_3222_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3222_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3221_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv919_3223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3226_inst
    process(conv919_3223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv919_3223(31 downto 0);
      type_cast_3226_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3228_inst
    process(conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv902_3097(31 downto 0);
      type_cast_3228_wire <= tmp_var; -- 
    end process;
    type_cast_3243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3243_inst_req_0;
      type_cast_3243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3243_inst_req_1;
      type_cast_3243_inst_ack_1<= rack(0);
      type_cast_3243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp927_3240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv928_3244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3258_inst
    process(conv919_3223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv919_3223(31 downto 0);
      type_cast_3258_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3260_inst
    process(add932_3255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add932_3255(31 downto 0);
      type_cast_3260_wire <= tmp_var; -- 
    end process;
    type_cast_3273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3273_inst_req_0;
      type_cast_3273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3273_inst_req_1;
      type_cast_3273_inst_ack_1<= rack(0);
      type_cast_3273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3272_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv939_3274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3278_inst_req_0;
      type_cast_3278_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3278_inst_req_1;
      type_cast_3278_inst_ack_1<= rack(0);
      type_cast_3278_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3277_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv943_3279,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3302_inst
    process(add951_3299) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add951_3299(31 downto 0);
      type_cast_3302_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3307_inst
    process(ASHR_i32_i32_3306_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3306_wire(31 downto 0);
      shr953_3308 <= tmp_var; -- 
    end process;
    type_cast_3312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3312_inst_req_0;
      type_cast_3312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3312_inst_req_1;
      type_cast_3312_inst_ack_1<= rack(0);
      type_cast_3312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3311_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom954_3313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3331_inst_req_0;
      type_cast_3331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3331_inst_req_1;
      type_cast_3331_inst_ack_1<= rack(0);
      type_cast_3331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3330_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv960_3332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3385_inst
    process(add978_3362) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add978_3362(31 downto 0);
      type_cast_3385_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3390_inst
    process(ASHR_i32_i32_3389_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3389_wire(31 downto 0);
      shr996_3391 <= tmp_var; -- 
    end process;
    type_cast_3395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3395_inst_req_0;
      type_cast_3395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3395_inst_req_1;
      type_cast_3395_inst_ack_1<= rack(0);
      type_cast_3395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3394_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom997_3396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3410_inst
    process(add994_3382) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add994_3382(31 downto 0);
      type_cast_3410_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3415_inst
    process(ASHR_i32_i32_3414_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3414_wire(31 downto 0);
      shr1001_3416 <= tmp_var; -- 
    end process;
    type_cast_3420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3420_inst_req_0;
      type_cast_3420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3420_inst_req_1;
      type_cast_3420_inst_ack_1<= rack(0);
      type_cast_3420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3419_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1002_3421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3438_inst_req_0;
      type_cast_3438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3438_inst_req_1;
      type_cast_3438_inst_ack_1<= rack(0);
      type_cast_3438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3437_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1008_3439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3448_inst
    process(add1009_3445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1009_3445(31 downto 0);
      type_cast_3448_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3450_inst
    process(conv880_3054) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv880_3054(31 downto 0);
      type_cast_3450_wire <= tmp_var; -- 
    end process;
    type_cast_3477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3477_inst_req_0;
      type_cast_3477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3477_inst_req_1;
      type_cast_3477_inst_ack_1<= rack(0);
      type_cast_3477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3476_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1023_3478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3484_inst_req_0;
      type_cast_3484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3484_inst_req_1;
      type_cast_3484_inst_ack_1<= rack(0);
      type_cast_3484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1024_3481,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1025_3485,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3504_inst_req_0;
      type_cast_3504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3504_inst_req_1;
      type_cast_3504_inst_ack_1<= rack(0);
      type_cast_3504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1031_3501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1036_3505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3521_inst_req_0;
      type_cast_3521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3521_inst_req_1;
      type_cast_3521_inst_ack_1<= rack(0);
      type_cast_3521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3520_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1039_3522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3528_inst_req_0;
      type_cast_3528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3528_inst_req_1;
      type_cast_3528_inst_ack_1<= rack(0);
      type_cast_3528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1040_3525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1041_3529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3562_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3562_inst_req_0;
      type_cast_3562_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3562_inst_req_1;
      type_cast_3562_inst_ack_1<= rack(0);
      type_cast_3562_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3562_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1017_3465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3562_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3569_inst_req_0;
      type_cast_3569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3569_inst_req_1;
      type_cast_3569_inst_ack_1<= rack(0);
      type_cast_3569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i844x_x2_3148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3569_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3571_inst_req_0;
      type_cast_3571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3571_inst_req_1;
      type_cast_3571_inst_ack_1<= rack(0);
      type_cast_3571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1036x_xi844x_x2_3510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3571_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3575_inst_req_0;
      type_cast_3575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3575_inst_req_1;
      type_cast_3575_inst_ack_1<= rack(0);
      type_cast_3575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j894x_x2_3517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3575_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3577_inst_req_0;
      type_cast_3577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3577_inst_req_1;
      type_cast_3577_inst_ack_1<= rack(0);
      type_cast_3577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j894x_x1_3154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3577_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3587_inst_req_0;
      type_cast_3587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3587_inst_req_1;
      type_cast_3587_inst_ack_1<= rack(0);
      type_cast_3587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1063_3584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1064_3588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3600_inst_req_0;
      type_cast_3600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3600_inst_req_1;
      type_cast_3600_inst_ack_1<= rack(0);
      type_cast_3600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1069_3597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1070_3601,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3640_inst_req_0;
      type_cast_3640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3640_inst_req_1;
      type_cast_3640_inst_ack_1<= rack(0);
      type_cast_3640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1079_3613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1104_3641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3644_inst_req_0;
      type_cast_3644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3644_inst_req_1;
      type_cast_3644_inst_ack_1<= rack(0);
      type_cast_3644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1063_3584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1106_3645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3654_inst
    process(sext1774_3651) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1774_3651(31 downto 0);
      type_cast_3654_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3659_inst
    process(ASHR_i32_i32_3658_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3658_wire(31 downto 0);
      conv1112_3660 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3669_inst
    process(sext1726_3666) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1726_3666(31 downto 0);
      type_cast_3669_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3674_inst
    process(ASHR_i32_i32_3673_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3673_wire(31 downto 0);
      conv1114_3675 <= tmp_var; -- 
    end process;
    type_cast_3683_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3683_inst_req_0;
      type_cast_3683_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3683_inst_req_1;
      type_cast_3683_inst_ack_1<= rack(0);
      type_cast_3683_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3683_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1075_3610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1126_3684,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3693_inst
    process(sext1775_3690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1775_3690(31 downto 0);
      type_cast_3693_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3698_inst
    process(ASHR_i32_i32_3697_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3697_wire(31 downto 0);
      conv1170_3699 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3719_inst
    process(sext1727_3716) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1727_3716(31 downto 0);
      type_cast_3719_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3724_inst
    process(ASHR_i32_i32_3723_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3723_wire(31 downto 0);
      conv1194_3725 <= tmp_var; -- 
    end process;
    type_cast_3731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3731_inst_req_0;
      type_cast_3731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3731_inst_req_1;
      type_cast_3731_inst_ack_1<= rack(0);
      type_cast_3731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1060x_x0x_xph_4132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3731_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3738_inst_req_0;
      type_cast_3738_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3738_inst_req_1;
      type_cast_3738_inst_ack_1<= rack(0);
      type_cast_3738_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3738_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1071_3607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3738_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3740_inst_req_0;
      type_cast_3740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3740_inst_req_1;
      type_cast_3740_inst_ack_1<= rack(0);
      type_cast_3740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1068x_x1x_xph_4139,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3740_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3744_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3744_inst_req_0;
      type_cast_3744_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3744_inst_req_1;
      type_cast_3744_inst_ack_1<= rack(0);
      type_cast_3744_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3744_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1118x_x0x_xph_4145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3744_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3746_inst_req_0;
      type_cast_3746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3746_inst_req_1;
      type_cast_3746_inst_ack_1<= rack(0);
      type_cast_3746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1065_3594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3746_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3751_inst_req_0;
      type_cast_3751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3751_inst_req_1;
      type_cast_3751_inst_ack_1<= rack(0);
      type_cast_3751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3750_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1124_3752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3755_inst
    process(conv1124_3752) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1124_3752(31 downto 0);
      type_cast_3755_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3757_inst
    process(conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1126_3684(31 downto 0);
      type_cast_3757_wire <= tmp_var; -- 
    end process;
    type_cast_3772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3772_inst_req_0;
      type_cast_3772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3772_inst_req_1;
      type_cast_3772_inst_ack_1<= rack(0);
      type_cast_3772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1132_3769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1133_3773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3793_inst
    process(conv1124_3752) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1124_3752(31 downto 0);
      type_cast_3793_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3795_inst
    process(add1138_3790) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1138_3790(31 downto 0);
      type_cast_3795_wire <= tmp_var; -- 
    end process;
    type_cast_3808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3808_inst_req_0;
      type_cast_3808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3808_inst_req_1;
      type_cast_3808_inst_ack_1<= rack(0);
      type_cast_3808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3807_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1143_3809,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3812_inst
    process(conv1143_3809) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1143_3809(31 downto 0);
      type_cast_3812_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3814_inst
    process(conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1126_3684(31 downto 0);
      type_cast_3814_wire <= tmp_var; -- 
    end process;
    type_cast_3829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3829_inst_req_0;
      type_cast_3829_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3829_inst_req_1;
      type_cast_3829_inst_ack_1<= rack(0);
      type_cast_3829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3829_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1151_3826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1152_3830,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3838_inst
    process(conv1143_3809) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1143_3809(31 downto 0);
      type_cast_3838_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3840_inst
    process(add1155_3835) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1155_3835(31 downto 0);
      type_cast_3840_wire <= tmp_var; -- 
    end process;
    type_cast_3853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3853_inst_req_0;
      type_cast_3853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3853_inst_req_1;
      type_cast_3853_inst_ack_1<= rack(0);
      type_cast_3853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3852_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1162_3854,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3858_inst_req_0;
      type_cast_3858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3858_inst_req_1;
      type_cast_3858_inst_ack_1<= rack(0);
      type_cast_3858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3857_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1166_3859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3882_inst
    process(add1174_3879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1174_3879(31 downto 0);
      type_cast_3882_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3887_inst
    process(ASHR_i32_i32_3886_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3886_wire(31 downto 0);
      shr1176_3888 <= tmp_var; -- 
    end process;
    type_cast_3892_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3892_inst_req_0;
      type_cast_3892_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3892_inst_req_1;
      type_cast_3892_inst_ack_1<= rack(0);
      type_cast_3892_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3892_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3891_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1177_3893,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3911_inst_req_0;
      type_cast_3911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3911_inst_req_1;
      type_cast_3911_inst_ack_1<= rack(0);
      type_cast_3911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3910_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1183_3912,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3965_inst
    process(add1201_3942) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1201_3942(31 downto 0);
      type_cast_3965_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3970_inst
    process(ASHR_i32_i32_3969_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3969_wire(31 downto 0);
      shr1219_3971 <= tmp_var; -- 
    end process;
    type_cast_3975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3975_inst_req_0;
      type_cast_3975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3975_inst_req_1;
      type_cast_3975_inst_ack_1<= rack(0);
      type_cast_3975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3974_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1220_3976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3990_inst
    process(add1217_3962) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1217_3962(31 downto 0);
      type_cast_3990_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3995_inst
    process(ASHR_i32_i32_3994_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3994_wire(31 downto 0);
      shr1224_3996 <= tmp_var; -- 
    end process;
    type_cast_4000_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4000_inst_req_0;
      type_cast_4000_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4000_inst_req_1;
      type_cast_4000_inst_ack_1<= rack(0);
      type_cast_4000_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4000_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3999_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1225_4001,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4018_inst_req_0;
      type_cast_4018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4018_inst_req_1;
      type_cast_4018_inst_ack_1<= rack(0);
      type_cast_4018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4017_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1231_4019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4028_inst
    process(add1232_4025) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1232_4025(31 downto 0);
      type_cast_4028_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4030_inst
    process(conv1104_3641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1104_3641(31 downto 0);
      type_cast_4030_wire <= tmp_var; -- 
    end process;
    type_cast_4057_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4057_inst_req_0;
      type_cast_4057_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4057_inst_req_1;
      type_cast_4057_inst_ack_1<= rack(0);
      type_cast_4057_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4057_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4056_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1246_4058,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4064_inst_req_0;
      type_cast_4064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4064_inst_req_1;
      type_cast_4064_inst_ack_1<= rack(0);
      type_cast_4064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1247_4061,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1248_4065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4078_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4078_inst_req_0;
      type_cast_4078_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4078_inst_req_1;
      type_cast_4078_inst_ack_1<= rack(0);
      type_cast_4078_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4078_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1253_4075,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1258_4079,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4094_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4094_inst_req_0;
      type_cast_4094_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4094_inst_req_1;
      type_cast_4094_inst_ack_1<= rack(0);
      type_cast_4094_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4094_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4093_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1261_4095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4101_inst_req_0;
      type_cast_4101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4101_inst_req_1;
      type_cast_4101_inst_ack_1<= rack(0);
      type_cast_4101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1262_4098,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1263_4102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4135_inst_req_0;
      type_cast_4135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4135_inst_req_1;
      type_cast_4135_inst_ack_1<= rack(0);
      type_cast_4135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1240_4045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4135_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4142_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4142_inst_req_0;
      type_cast_4142_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4142_inst_req_1;
      type_cast_4142_inst_ack_1<= rack(0);
      type_cast_4142_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4142_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1068x_x2_3735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4142_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4144_inst_req_0;
      type_cast_4144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4144_inst_req_1;
      type_cast_4144_inst_ack_1<= rack(0);
      type_cast_4144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1258x_xi1068x_x2_4084,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4144_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4148_inst_req_0;
      type_cast_4148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4148_inst_req_1;
      type_cast_4148_inst_ack_1<= rack(0);
      type_cast_4148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1118x_x1_3741,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4148_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4150_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4150_inst_req_0;
      type_cast_4150_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4150_inst_req_1;
      type_cast_4150_inst_ack_1<= rack(0);
      type_cast_4150_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4150_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1118x_x2_4090,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4150_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4160_inst_req_0;
      type_cast_4160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4160_inst_req_1;
      type_cast_4160_inst_ack_1<= rack(0);
      type_cast_4160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1287_4157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1288_4161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4209_inst_req_0;
      type_cast_4209_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4209_inst_req_1;
      type_cast_4209_inst_ack_1<= rack(0);
      type_cast_4209_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1298_4179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1323_4210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4213_inst_req_0;
      type_cast_4213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4213_inst_req_1;
      type_cast_4213_inst_ack_1<= rack(0);
      type_cast_4213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1302_4182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1325_4214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4223_inst
    process(sext1776_4220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1776_4220(31 downto 0);
      type_cast_4223_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4228_inst
    process(ASHR_i32_i32_4227_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4227_wire(31 downto 0);
      conv1331_4229 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4238_inst
    process(sext1728_4235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1728_4235(31 downto 0);
      type_cast_4238_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4243_inst
    process(ASHR_i32_i32_4242_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4242_wire(31 downto 0);
      conv1333_4244 <= tmp_var; -- 
    end process;
    type_cast_4252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4252_inst_req_0;
      type_cast_4252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4252_inst_req_1;
      type_cast_4252_inst_ack_1<= rack(0);
      type_cast_4252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1294_4176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1345_4253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4262_inst
    process(sext1777_4259) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1777_4259(31 downto 0);
      type_cast_4262_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4267_inst
    process(ASHR_i32_i32_4266_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4266_wire(31 downto 0);
      conv1388_4268 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4288_inst
    process(sext1729_4285) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1729_4285(31 downto 0);
      type_cast_4288_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4293_inst
    process(ASHR_i32_i32_4292_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4292_wire(31 downto 0);
      conv1412_4294 <= tmp_var; -- 
    end process;
    type_cast_4303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4303_inst_req_0;
      type_cast_4303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4303_inst_req_1;
      type_cast_4303_inst_ack_1<= rack(0);
      type_cast_4303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1282x_x0x_xph_4691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4303_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4307_inst_req_0;
      type_cast_4307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4307_inst_req_1;
      type_cast_4307_inst_ack_1<= rack(0);
      type_cast_4307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul1290_4173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4307_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4309_inst_req_0;
      type_cast_4309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4309_inst_req_1;
      type_cast_4309_inst_ack_1<= rack(0);
      type_cast_4309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1286x_x1x_xph_4698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4316_inst_req_0;
      type_cast_4316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4316_inst_req_1;
      type_cast_4316_inst_ack_1<= rack(0);
      type_cast_4316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1337x_x0x_xph_4704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4316_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4321_inst_req_0;
      type_cast_4321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4321_inst_req_1;
      type_cast_4321_inst_ack_1<= rack(0);
      type_cast_4321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4320_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1343_4322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4325_inst
    process(conv1343_4322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1343_4322(31 downto 0);
      type_cast_4325_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4327_inst
    process(conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1345_4253(31 downto 0);
      type_cast_4327_wire <= tmp_var; -- 
    end process;
    type_cast_4342_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4342_inst_req_0;
      type_cast_4342_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4342_inst_req_1;
      type_cast_4342_inst_ack_1<= rack(0);
      type_cast_4342_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4342_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1351_4339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1352_4343,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4351_inst
    process(conv1343_4322) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1343_4322(31 downto 0);
      type_cast_4351_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4353_inst
    process(add1355_4348) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1355_4348(31 downto 0);
      type_cast_4353_wire <= tmp_var; -- 
    end process;
    type_cast_4366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4366_inst_req_0;
      type_cast_4366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4366_inst_req_1;
      type_cast_4366_inst_ack_1<= rack(0);
      type_cast_4366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4365_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1360_4367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4370_inst
    process(conv1360_4367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1360_4367(31 downto 0);
      type_cast_4370_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4372_inst
    process(conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1345_4253(31 downto 0);
      type_cast_4372_wire <= tmp_var; -- 
    end process;
    type_cast_4387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4387_inst_req_0;
      type_cast_4387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4387_inst_req_1;
      type_cast_4387_inst_ack_1<= rack(0);
      type_cast_4387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1368_4384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1369_4388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4402_inst
    process(conv1360_4367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1360_4367(31 downto 0);
      type_cast_4402_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4404_inst
    process(add1373_4399) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1373_4399(31 downto 0);
      type_cast_4404_wire <= tmp_var; -- 
    end process;
    type_cast_4417_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4417_inst_req_0;
      type_cast_4417_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4417_inst_req_1;
      type_cast_4417_inst_ack_1<= rack(0);
      type_cast_4417_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4417_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4416_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1380_4418,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4422_inst_req_0;
      type_cast_4422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4422_inst_req_1;
      type_cast_4422_inst_ack_1<= rack(0);
      type_cast_4422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4421_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1384_4423,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4446_inst
    process(add1392_4443) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1392_4443(31 downto 0);
      type_cast_4446_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4451_inst
    process(ASHR_i32_i32_4450_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4450_wire(31 downto 0);
      shr1394_4452 <= tmp_var; -- 
    end process;
    type_cast_4456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4456_inst_req_0;
      type_cast_4456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4456_inst_req_1;
      type_cast_4456_inst_ack_1<= rack(0);
      type_cast_4456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4455_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1395_4457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4475_inst_req_0;
      type_cast_4475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4475_inst_req_1;
      type_cast_4475_inst_ack_1<= rack(0);
      type_cast_4475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4474_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1401_4476,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4529_inst
    process(add1419_4506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1419_4506(31 downto 0);
      type_cast_4529_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4534_inst
    process(ASHR_i32_i32_4533_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4533_wire(31 downto 0);
      shr1437_4535 <= tmp_var; -- 
    end process;
    type_cast_4539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4539_inst_req_0;
      type_cast_4539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4539_inst_req_1;
      type_cast_4539_inst_ack_1<= rack(0);
      type_cast_4539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4538_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1438_4540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4554_inst
    process(add1435_4526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1435_4526(31 downto 0);
      type_cast_4554_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4559_inst
    process(ASHR_i32_i32_4558_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4558_wire(31 downto 0);
      shr1442_4560 <= tmp_var; -- 
    end process;
    type_cast_4564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4564_inst_req_0;
      type_cast_4564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4564_inst_req_1;
      type_cast_4564_inst_ack_1<= rack(0);
      type_cast_4564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4563_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1443_4565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4582_inst_req_0;
      type_cast_4582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4582_inst_req_1;
      type_cast_4582_inst_ack_1<= rack(0);
      type_cast_4582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4581_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1449_4583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4592_inst
    process(add1450_4589) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1450_4589(31 downto 0);
      type_cast_4592_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4594_inst
    process(conv1323_4210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1323_4210(31 downto 0);
      type_cast_4594_wire <= tmp_var; -- 
    end process;
    type_cast_4621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4621_inst_req_0;
      type_cast_4621_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4621_inst_req_1;
      type_cast_4621_inst_ack_1<= rack(0);
      type_cast_4621_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4621_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4620_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1464_4622,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4628_inst_req_0;
      type_cast_4628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4628_inst_req_1;
      type_cast_4628_inst_ack_1<= rack(0);
      type_cast_4628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4628_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1465_4625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1466_4629,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4648_inst_req_0;
      type_cast_4648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4648_inst_req_1;
      type_cast_4648_inst_ack_1<= rack(0);
      type_cast_4648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1472_4645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1477_4649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4665_inst_req_0;
      type_cast_4665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4665_inst_req_1;
      type_cast_4665_inst_ack_1<= rack(0);
      type_cast_4665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4664_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1480_4666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4672_inst_req_0;
      type_cast_4672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4672_inst_req_1;
      type_cast_4672_inst_ack_1<= rack(0);
      type_cast_4672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1481_4669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1482_4673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4694_inst_req_0;
      type_cast_4694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4694_inst_req_1;
      type_cast_4694_inst_ack_1<= rack(0);
      type_cast_4694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1458_4609,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4694_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4701_inst_req_0;
      type_cast_4701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4701_inst_req_1;
      type_cast_4701_inst_ack_1<= rack(0);
      type_cast_4701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1286x_x2_4304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4701_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4703_inst_req_0;
      type_cast_4703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4703_inst_req_1;
      type_cast_4703_inst_ack_1<= rack(0);
      type_cast_4703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1477x_xi1286x_x2_4654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4703_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4707_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4707_inst_req_0;
      type_cast_4707_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4707_inst_req_1;
      type_cast_4707_inst_ack_1<= rack(0);
      type_cast_4707_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4707_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1337x_x1_4310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4707_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4709_inst_req_0;
      type_cast_4709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4709_inst_req_1;
      type_cast_4709_inst_ack_1<= rack(0);
      type_cast_4709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1337x_x2_4661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4709_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4719_inst_req_0;
      type_cast_4719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4719_inst_req_1;
      type_cast_4719_inst_ack_1<= rack(0);
      type_cast_4719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1502_4716,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1503_4720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4732_inst_req_0;
      type_cast_4732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4732_inst_req_1;
      type_cast_4732_inst_ack_1<= rack(0);
      type_cast_4732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1508_4729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1509_4733,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4778_inst_req_0;
      type_cast_4778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4778_inst_req_1;
      type_cast_4778_inst_ack_1<= rack(0);
      type_cast_4778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1519_4751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1544_4779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4782_inst_req_0;
      type_cast_4782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4782_inst_req_1;
      type_cast_4782_inst_ack_1<= rack(0);
      type_cast_4782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1502_4716,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1546_4783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4792_inst
    process(sext1778_4789) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1778_4789(31 downto 0);
      type_cast_4792_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4797_inst
    process(ASHR_i32_i32_4796_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4796_wire(31 downto 0);
      conv1552_4798 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4807_inst
    process(sext1730_4804) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1730_4804(31 downto 0);
      type_cast_4807_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4812_inst
    process(ASHR_i32_i32_4811_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4811_wire(31 downto 0);
      conv1554_4813 <= tmp_var; -- 
    end process;
    type_cast_4821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4821_inst_req_0;
      type_cast_4821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4821_inst_req_1;
      type_cast_4821_inst_ack_1<= rack(0);
      type_cast_4821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1515_4748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1566_4822,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4831_inst
    process(sext1779_4828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1779_4828(31 downto 0);
      type_cast_4831_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4836_inst
    process(ASHR_i32_i32_4835_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4835_wire(31 downto 0);
      conv1608_4837 <= tmp_var; -- 
    end process;
    -- interlock type_cast_4857_inst
    process(sext1731_4854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1731_4854(31 downto 0);
      type_cast_4857_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4862_inst
    process(ASHR_i32_i32_4861_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_4861_wire(31 downto 0);
      conv1632_4863 <= tmp_var; -- 
    end process;
    type_cast_4872_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4872_inst_req_0;
      type_cast_4872_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4872_inst_req_1;
      type_cast_4872_inst_ack_1<= rack(0);
      type_cast_4872_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4872_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1499x_x0x_xph_5246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4872_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4876_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4876_inst_req_0;
      type_cast_4876_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4876_inst_req_1;
      type_cast_4876_inst_ack_1<= rack(0);
      type_cast_4876_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4876_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1507x_x1x_xph_5253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4876_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4878_inst_req_0;
      type_cast_4878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4878_inst_req_1;
      type_cast_4878_inst_ack_1<= rack(0);
      type_cast_4878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4878_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1511_4745,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4878_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4882_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4882_inst_req_0;
      type_cast_4882_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4882_inst_req_1;
      type_cast_4882_inst_ack_1<= rack(0);
      type_cast_4882_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4882_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1504_4726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4882_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4884_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4884_inst_req_0;
      type_cast_4884_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4884_inst_req_1;
      type_cast_4884_inst_ack_1<= rack(0);
      type_cast_4884_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4884_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1558x_x0x_xph_5259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_4884_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4889_inst_req_0;
      type_cast_4889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4889_inst_req_1;
      type_cast_4889_inst_ack_1<= rack(0);
      type_cast_4889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4888_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1564_4890,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4893_inst
    process(conv1564_4890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1564_4890(31 downto 0);
      type_cast_4893_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4895_inst
    process(conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1566_4822(31 downto 0);
      type_cast_4895_wire <= tmp_var; -- 
    end process;
    type_cast_4910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4910_inst_req_0;
      type_cast_4910_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4910_inst_req_1;
      type_cast_4910_inst_ack_1<= rack(0);
      type_cast_4910_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4910_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1572_4907,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1573_4911,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4919_inst
    process(conv1564_4890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1564_4890(31 downto 0);
      type_cast_4919_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4921_inst
    process(add1576_4916) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1576_4916(31 downto 0);
      type_cast_4921_wire <= tmp_var; -- 
    end process;
    type_cast_4934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4934_inst_req_0;
      type_cast_4934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4934_inst_req_1;
      type_cast_4934_inst_ack_1<= rack(0);
      type_cast_4934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4933_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1581_4935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4938_inst
    process(conv1581_4935) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1581_4935(31 downto 0);
      type_cast_4938_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4940_inst
    process(conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1566_4822(31 downto 0);
      type_cast_4940_wire <= tmp_var; -- 
    end process;
    type_cast_4955_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4955_inst_req_0;
      type_cast_4955_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4955_inst_req_1;
      type_cast_4955_inst_ack_1<= rack(0);
      type_cast_4955_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4955_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1589_4952,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1590_4956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_4964_inst
    process(conv1581_4935) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1581_4935(31 downto 0);
      type_cast_4964_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_4966_inst
    process(add1593_4961) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1593_4961(31 downto 0);
      type_cast_4966_wire <= tmp_var; -- 
    end process;
    type_cast_4979_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4979_inst_req_0;
      type_cast_4979_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4979_inst_req_1;
      type_cast_4979_inst_ack_1<= rack(0);
      type_cast_4979_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4979_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4978_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1600_4980,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_4984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_4984_inst_req_0;
      type_cast_4984_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_4984_inst_req_1;
      type_cast_4984_inst_ack_1<= rack(0);
      type_cast_4984_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_4984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_4983_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1604_4985,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5008_inst
    process(add1612_5005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1612_5005(31 downto 0);
      type_cast_5008_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5013_inst
    process(ASHR_i32_i32_5012_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_5012_wire(31 downto 0);
      shr1614_5014 <= tmp_var; -- 
    end process;
    type_cast_5018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5018_inst_req_0;
      type_cast_5018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5018_inst_req_1;
      type_cast_5018_inst_ack_1<= rack(0);
      type_cast_5018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5017_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1615_5019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5037_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5037_inst_req_0;
      type_cast_5037_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5037_inst_req_1;
      type_cast_5037_inst_ack_1<= rack(0);
      type_cast_5037_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5037_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5036_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1621_5038,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5091_inst
    process(add1639_5068) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1639_5068(31 downto 0);
      type_cast_5091_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5096_inst
    process(ASHR_i32_i32_5095_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_5095_wire(31 downto 0);
      shr1657_5097 <= tmp_var; -- 
    end process;
    type_cast_5101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5101_inst_req_0;
      type_cast_5101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5101_inst_req_1;
      type_cast_5101_inst_ack_1<= rack(0);
      type_cast_5101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5100_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1658_5102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5116_inst
    process(add1655_5088) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1655_5088(31 downto 0);
      type_cast_5116_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5121_inst
    process(ASHR_i32_i32_5120_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_5120_wire(31 downto 0);
      shr1662_5122 <= tmp_var; -- 
    end process;
    type_cast_5126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5126_inst_req_0;
      type_cast_5126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5126_inst_req_1;
      type_cast_5126_inst_ack_1<= rack(0);
      type_cast_5126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5125_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1663_5127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5144_inst_req_0;
      type_cast_5144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5144_inst_req_1;
      type_cast_5144_inst_ack_1<= rack(0);
      type_cast_5144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5143_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1669_5145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_5154_inst
    process(add1670_5151) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1670_5151(31 downto 0);
      type_cast_5154_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_5156_inst
    process(conv1544_4779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1544_4779(31 downto 0);
      type_cast_5156_wire <= tmp_var; -- 
    end process;
    type_cast_5183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5183_inst_req_0;
      type_cast_5183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5183_inst_req_1;
      type_cast_5183_inst_ack_1<= rack(0);
      type_cast_5183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5182_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1684_5184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5190_inst_req_0;
      type_cast_5190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5190_inst_req_1;
      type_cast_5190_inst_ack_1<= rack(0);
      type_cast_5190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1685_5187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1686_5191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5204_inst_req_0;
      type_cast_5204_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5204_inst_req_1;
      type_cast_5204_inst_ack_1<= rack(0);
      type_cast_5204_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1691_5201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1696_5205,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5220_inst_req_0;
      type_cast_5220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5220_inst_req_1;
      type_cast_5220_inst_ack_1<= rack(0);
      type_cast_5220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_5219_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1699_5221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5227_inst_req_0;
      type_cast_5227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5227_inst_req_1;
      type_cast_5227_inst_ack_1<= rack(0);
      type_cast_5227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1700_5224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1701_5228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5252_inst_req_0;
      type_cast_5252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5252_inst_req_1;
      type_cast_5252_inst_ack_1<= rack(0);
      type_cast_5252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1678_5171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5252_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5256_inst_req_0;
      type_cast_5256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5256_inst_req_1;
      type_cast_5256_inst_ack_1<= rack(0);
      type_cast_5256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1507x_x2_4873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5256_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5258_inst_req_0;
      type_cast_5258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5258_inst_req_1;
      type_cast_5258_inst_ack_1<= rack(0);
      type_cast_5258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1696x_xi1507x_x2_5210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5258_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5262_inst_req_0;
      type_cast_5262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5262_inst_req_1;
      type_cast_5262_inst_ack_1<= rack(0);
      type_cast_5262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1558x_x1_4879,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5262_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_5264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_5264_inst_req_0;
      type_cast_5264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_5264_inst_req_1;
      type_cast_5264_inst_ack_1<= rack(0);
      type_cast_5264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_5264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1558x_x2_5216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_5264_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_731_inst_req_0;
      type_cast_731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_731_inst_req_1;
      type_cast_731_inst_ack_1<= rack(0);
      type_cast_731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_769_inst_req_0;
      type_cast_769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_769_inst_req_1;
      type_cast_769_inst_ack_1<= rack(0);
      type_cast_769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_766,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_810_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_810_inst_req_0;
      type_cast_810_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_810_inst_req_1;
      type_cast_810_inst_ack_1<= rack(0);
      type_cast_810_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_810_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_811,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_814_inst_req_0;
      type_cast_814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_814_inst_req_1;
      type_cast_814_inst_ack_1<= rack(0);
      type_cast_814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp15_783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_825_inst
    process(sext1764_821) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1764_821(31 downto 0);
      type_cast_825_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_830_inst
    process(ASHR_i32_i32_829_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_829_wire(31 downto 0);
      conv37_831 <= tmp_var; -- 
    end process;
    -- interlock type_cast_840_inst
    process(sext_837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_837(31 downto 0);
      type_cast_840_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_845_inst
    process(ASHR_i32_i32_844_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_844_wire(31 downto 0);
      conv39_846 <= tmp_var; -- 
    end process;
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_864_inst
    process(sext1765_861) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1765_861(31 downto 0);
      type_cast_864_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_869_inst
    process(ASHR_i32_i32_868_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_868_wire(31 downto 0);
      conv86_870 <= tmp_var; -- 
    end process;
    -- interlock type_cast_890_inst
    process(sext1717_887) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1717_887(31 downto 0);
      type_cast_890_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_895_inst
    process(ASHR_i32_i32_894_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_894_wire(31 downto 0);
      conv104_896 <= tmp_var; -- 
    end process;
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_905_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_912_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_912_inst_req_0;
      type_cast_912_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_912_inst_req_1;
      type_cast_912_inst_ack_1<= rack(0);
      type_cast_912_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_912_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1x_xph_1313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_912_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_919_inst_req_0;
      type_cast_919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_919_inst_req_1;
      type_cast_919_inst_ack_1<= rack(0);
      type_cast_919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_1319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_919_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_924_inst_req_0;
      type_cast_924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_924_inst_req_1;
      type_cast_924_inst_ack_1<= rack(0);
      type_cast_924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_923_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_928_inst
    process(conv46_925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_925(31 downto 0);
      type_cast_928_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_930_inst
    process(conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_855(31 downto 0);
      type_cast_930_wire <= tmp_var; -- 
    end process;
    type_cast_945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_945_inst_req_0;
      type_cast_945_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_945_inst_req_1;
      type_cast_945_inst_ack_1<= rack(0);
      type_cast_945_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp52_942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_946,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_960_inst
    process(conv46_925) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv46_925(31 downto 0);
      type_cast_960_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_962_inst
    process(add_957) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_957(31 downto 0);
      type_cast_962_wire <= tmp_var; -- 
    end process;
    type_cast_975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_975_inst_req_0;
      type_cast_975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_975_inst_req_1;
      type_cast_975_inst_ack_1<= rack(0);
      type_cast_975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_974_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_979_inst
    process(conv60_976) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv60_976(31 downto 0);
      type_cast_979_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_981_inst
    process(conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv48_855(31 downto 0);
      type_cast_981_wire <= tmp_var; -- 
    end process;
    type_cast_996_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_996_inst_req_0;
      type_cast_996_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_996_inst_req_1;
      type_cast_996_inst_ack_1<= rack(0);
      type_cast_996_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_996_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp68_993,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_997,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_col_high_1234_gather_scatter
    process(LOAD_col_high_1234_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1234_data_0;
      ov(7 downto 0) := iv;
      tmp154_1235 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1331_gather_scatter
    process(LOAD_col_high_1331_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1331_data_0;
      ov(7 downto 0) := iv;
      tmp189_1332 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1555_gather_scatter
    process(LOAD_col_high_1555_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1555_data_0;
      ov(7 downto 0) := iv;
      tmp272_1556 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1790_gather_scatter
    process(LOAD_col_high_1790_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1790_data_0;
      ov(7 downto 0) := iv;
      tmp368_1791 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_1899_gather_scatter
    process(LOAD_col_high_1899_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_1899_data_0;
      ov(7 downto 0) := iv;
      tmp421_1900 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2107_gather_scatter
    process(LOAD_col_high_2107_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2107_data_0;
      ov(7 downto 0) := iv;
      tmp488_2108 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2348_gather_scatter
    process(LOAD_col_high_2348_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2348_data_0;
      ov(7 downto 0) := iv;
      tmp585_2349 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2445_gather_scatter
    process(LOAD_col_high_2445_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2445_data_0;
      ov(7 downto 0) := iv;
      tmp623_2446 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2681_gather_scatter
    process(LOAD_col_high_2681_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2681_data_0;
      ov(7 downto 0) := iv;
      tmp710_2682 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_2916_gather_scatter
    process(LOAD_col_high_2916_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_2916_data_0;
      ov(7 downto 0) := iv;
      tmp806_2917 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3025_gather_scatter
    process(LOAD_col_high_3025_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3025_data_0;
      ov(7 downto 0) := iv;
      tmp859_3026 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3239_gather_scatter
    process(LOAD_col_high_3239_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3239_data_0;
      ov(7 downto 0) := iv;
      tmp927_3240 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3480_gather_scatter
    process(LOAD_col_high_3480_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3480_data_0;
      ov(7 downto 0) := iv;
      tmp1024_3481 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3583_gather_scatter
    process(LOAD_col_high_3583_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3583_data_0;
      ov(7 downto 0) := iv;
      tmp1063_3584 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_3825_gather_scatter
    process(LOAD_col_high_3825_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_3825_data_0;
      ov(7 downto 0) := iv;
      tmp1151_3826 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4060_gather_scatter
    process(LOAD_col_high_4060_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4060_data_0;
      ov(7 downto 0) := iv;
      tmp1247_4061 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4181_gather_scatter
    process(LOAD_col_high_4181_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4181_data_0;
      ov(7 downto 0) := iv;
      tmp1302_4182 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4383_gather_scatter
    process(LOAD_col_high_4383_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4383_data_0;
      ov(7 downto 0) := iv;
      tmp1368_4384 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4624_gather_scatter
    process(LOAD_col_high_4624_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4624_data_0;
      ov(7 downto 0) := iv;
      tmp1465_4625 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4715_gather_scatter
    process(LOAD_col_high_4715_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4715_data_0;
      ov(7 downto 0) := iv;
      tmp1502_4716 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_4951_gather_scatter
    process(LOAD_col_high_4951_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_4951_data_0;
      ov(7 downto 0) := iv;
      tmp1589_4952 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_5186_gather_scatter
    process(LOAD_col_high_5186_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_5186_data_0;
      ov(7 downto 0) := iv;
      tmp1685_5187 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_782_gather_scatter
    process(LOAD_col_high_782_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_782_data_0;
      ov(7 downto 0) := iv;
      tmp15_783 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_col_high_992_gather_scatter
    process(LOAD_col_high_992_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_col_high_992_data_0;
      ov(7 downto 0) := iv;
      tmp68_993 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_1347_gather_scatter
    process(LOAD_depth_high_1347_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_1347_data_0;
      ov(7 downto 0) := iv;
      tmp201_1348 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_1896_gather_scatter
    process(LOAD_depth_high_1896_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_1896_data_0;
      ov(7 downto 0) := iv;
      tmp417_1897 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_2474_gather_scatter
    process(LOAD_depth_high_2474_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_2474_data_0;
      ov(7 downto 0) := iv;
      tmp639_2475 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_3022_gather_scatter
    process(LOAD_depth_high_3022_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_3022_data_0;
      ov(7 downto 0) := iv;
      tmp855_3023 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_3612_gather_scatter
    process(LOAD_depth_high_3612_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_3612_data_0;
      ov(7 downto 0) := iv;
      tmp1079_3613 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_4178_gather_scatter
    process(LOAD_depth_high_4178_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_4178_data_0;
      ov(7 downto 0) := iv;
      tmp1298_4179 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_4750_gather_scatter
    process(LOAD_depth_high_4750_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_4750_data_0;
      ov(7 downto 0) := iv;
      tmp1519_4751 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_depth_high_779_gather_scatter
    process(LOAD_depth_high_779_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_depth_high_779_data_0;
      ov(7 downto 0) := iv;
      tmp12_780 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1344_gather_scatter
    process(LOAD_pad_1344_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1344_data_0;
      ov(7 downto 0) := iv;
      tmp197_1345 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1893_gather_scatter
    process(LOAD_pad_1893_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1893_data_0;
      ov(7 downto 0) := iv;
      tmp413_1894 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_2471_gather_scatter
    process(LOAD_pad_2471_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2471_data_0;
      ov(7 downto 0) := iv;
      tmp635_2472 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3019_gather_scatter
    process(LOAD_pad_3019_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3019_data_0;
      ov(7 downto 0) := iv;
      tmp851_3020 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3609_gather_scatter
    process(LOAD_pad_3609_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3609_data_0;
      ov(7 downto 0) := iv;
      tmp1075_3610 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_4175_gather_scatter
    process(LOAD_pad_4175_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_4175_data_0;
      ov(7 downto 0) := iv;
      tmp1294_4176 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_4747_gather_scatter
    process(LOAD_pad_4747_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_4747_data_0;
      ov(7 downto 0) := iv;
      tmp1515_4748 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_776_gather_scatter
    process(LOAD_pad_776_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_776_data_0;
      ov(7 downto 0) := iv;
      tmp9_777 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1278_gather_scatter
    process(LOAD_row_high_1278_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1278_data_0;
      ov(7 downto 0) := iv;
      tmp169_1279 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1504_gather_scatter
    process(LOAD_row_high_1504_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1504_data_0;
      ov(7 downto 0) := iv;
      tmp254_1505 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1827_gather_scatter
    process(LOAD_row_high_1827_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1827_data_0;
      ov(7 downto 0) := iv;
      tmp383_1828 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_1880_gather_scatter
    process(LOAD_row_high_1880_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_1880_data_0;
      ov(7 downto 0) := iv;
      tmp407_1881 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2056_gather_scatter
    process(LOAD_row_high_2056_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2056_data_0;
      ov(7 downto 0) := iv;
      tmp470_2057 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2392_gather_scatter
    process(LOAD_row_high_2392_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2392_data_0;
      ov(7 downto 0) := iv;
      tmp601_2393 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2458_gather_scatter
    process(LOAD_row_high_2458_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2458_data_0;
      ov(7 downto 0) := iv;
      tmp629_2459 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2630_gather_scatter
    process(LOAD_row_high_2630_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2630_data_0;
      ov(7 downto 0) := iv;
      tmp692_2631 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_2953_gather_scatter
    process(LOAD_row_high_2953_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_2953_data_0;
      ov(7 downto 0) := iv;
      tmp821_2954 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3006_gather_scatter
    process(LOAD_row_high_3006_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3006_data_0;
      ov(7 downto 0) := iv;
      tmp845_3007 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3182_gather_scatter
    process(LOAD_row_high_3182_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3182_data_0;
      ov(7 downto 0) := iv;
      tmp908_3183 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3524_gather_scatter
    process(LOAD_row_high_3524_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3524_data_0;
      ov(7 downto 0) := iv;
      tmp1040_3525 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3596_gather_scatter
    process(LOAD_row_high_3596_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3596_data_0;
      ov(7 downto 0) := iv;
      tmp1069_3597 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_3768_gather_scatter
    process(LOAD_row_high_3768_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_3768_data_0;
      ov(7 downto 0) := iv;
      tmp1132_3769 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4097_gather_scatter
    process(LOAD_row_high_4097_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4097_data_0;
      ov(7 downto 0) := iv;
      tmp1262_4098 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4156_gather_scatter
    process(LOAD_row_high_4156_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4156_data_0;
      ov(7 downto 0) := iv;
      tmp1287_4157 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4338_gather_scatter
    process(LOAD_row_high_4338_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4338_data_0;
      ov(7 downto 0) := iv;
      tmp1351_4339 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4668_gather_scatter
    process(LOAD_row_high_4668_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4668_data_0;
      ov(7 downto 0) := iv;
      tmp1481_4669 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4728_gather_scatter
    process(LOAD_row_high_4728_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4728_data_0;
      ov(7 downto 0) := iv;
      tmp1508_4729 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_4906_gather_scatter
    process(LOAD_row_high_4906_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_4906_data_0;
      ov(7 downto 0) := iv;
      tmp1572_4907 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_5223_gather_scatter
    process(LOAD_row_high_5223_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_5223_data_0;
      ov(7 downto 0) := iv;
      tmp1700_5224 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_row_high_941_gather_scatter
    process(LOAD_row_high_941_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_row_high_941_data_0;
      ov(7 downto 0) := iv;
      tmp52_942 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_col_high_752_gather_scatter
    process(conv2_751) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv2_751;
      ov(7 downto 0) := iv;
      STORE_col_high_752_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_depth_high_771_gather_scatter
    process(conv4_770) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4_770;
      ov(7 downto 0) := iv;
      STORE_depth_high_771_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_row_high_733_gather_scatter
    process(conv_732) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_732;
      ov(7 downto 0) := iv;
      STORE_row_high_733_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_index_1_rename
    process(R_idxprom_1071_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1071_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1071_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_index_1_resize
    process(idxprom_1067) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1067;
      ov := iv(13 downto 0);
      R_idxprom_1071_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_root_address_inst
    process(array_obj_ref_1072_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1072_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1072_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_index_1_rename
    process(R_idxprom130_1154_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom130_1154_resized;
      ov(13 downto 0) := iv;
      R_idxprom130_1154_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_index_1_resize
    process(idxprom130_1150) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom130_1150;
      ov := iv(13 downto 0);
      R_idxprom130_1154_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1155_root_address_inst
    process(array_obj_ref_1155_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1155_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1155_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1180_index_1_rename
    process(R_idxprom135_1179_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom135_1179_resized;
      ov(13 downto 0) := iv;
      R_idxprom135_1179_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1180_index_1_resize
    process(idxprom135_1175) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom135_1175;
      ov := iv(13 downto 0);
      R_idxprom135_1179_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1180_root_address_inst
    process(array_obj_ref_1180_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1180_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1180_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1628_index_1_rename
    process(R_idxprom298_1627_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom298_1627_resized;
      ov(13 downto 0) := iv;
      R_idxprom298_1627_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1628_index_1_resize
    process(idxprom298_1623) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom298_1623;
      ov := iv(13 downto 0);
      R_idxprom298_1627_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1628_root_address_inst
    process(array_obj_ref_1628_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1628_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1628_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1711_index_1_rename
    process(R_idxprom341_1710_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom341_1710_resized;
      ov(13 downto 0) := iv;
      R_idxprom341_1710_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1711_index_1_resize
    process(idxprom341_1706) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom341_1706;
      ov := iv(13 downto 0);
      R_idxprom341_1710_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1711_root_address_inst
    process(array_obj_ref_1711_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1711_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1711_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1736_index_1_rename
    process(R_idxprom346_1735_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom346_1735_resized;
      ov(13 downto 0) := iv;
      R_idxprom346_1735_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1736_index_1_resize
    process(idxprom346_1731) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom346_1731;
      ov := iv(13 downto 0);
      R_idxprom346_1735_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1736_root_address_inst
    process(array_obj_ref_1736_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1736_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1736_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2186_index_1_rename
    process(R_idxprom515_2185_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom515_2185_resized;
      ov(13 downto 0) := iv;
      R_idxprom515_2185_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2186_index_1_resize
    process(idxprom515_2181) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom515_2181;
      ov := iv(13 downto 0);
      R_idxprom515_2185_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2186_root_address_inst
    process(array_obj_ref_2186_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2186_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2186_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2269_index_1_rename
    process(R_idxprom558_2268_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom558_2268_resized;
      ov(13 downto 0) := iv;
      R_idxprom558_2268_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2269_index_1_resize
    process(idxprom558_2264) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom558_2264;
      ov := iv(13 downto 0);
      R_idxprom558_2268_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2269_root_address_inst
    process(array_obj_ref_2269_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2269_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2269_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2294_index_1_rename
    process(R_idxprom563_2293_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom563_2293_resized;
      ov(13 downto 0) := iv;
      R_idxprom563_2293_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2294_index_1_resize
    process(idxprom563_2289) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom563_2289;
      ov := iv(13 downto 0);
      R_idxprom563_2293_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2294_root_address_inst
    process(array_obj_ref_2294_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2294_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2294_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2754_index_1_rename
    process(R_idxprom736_2753_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom736_2753_resized;
      ov(13 downto 0) := iv;
      R_idxprom736_2753_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2754_index_1_resize
    process(idxprom736_2749) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom736_2749;
      ov := iv(13 downto 0);
      R_idxprom736_2753_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2754_root_address_inst
    process(array_obj_ref_2754_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2754_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2754_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2837_index_1_rename
    process(R_idxprom779_2836_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom779_2836_resized;
      ov(13 downto 0) := iv;
      R_idxprom779_2836_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2837_index_1_resize
    process(idxprom779_2832) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom779_2832;
      ov := iv(13 downto 0);
      R_idxprom779_2836_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2837_root_address_inst
    process(array_obj_ref_2837_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2837_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2837_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2862_index_1_rename
    process(R_idxprom784_2861_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom784_2861_resized;
      ov(13 downto 0) := iv;
      R_idxprom784_2861_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2862_index_1_resize
    process(idxprom784_2857) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom784_2857;
      ov := iv(13 downto 0);
      R_idxprom784_2861_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2862_root_address_inst
    process(array_obj_ref_2862_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2862_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2862_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3318_index_1_rename
    process(R_idxprom954_3317_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom954_3317_resized;
      ov(13 downto 0) := iv;
      R_idxprom954_3317_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3318_index_1_resize
    process(idxprom954_3313) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom954_3313;
      ov := iv(13 downto 0);
      R_idxprom954_3317_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3318_root_address_inst
    process(array_obj_ref_3318_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3318_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3318_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3401_index_1_rename
    process(R_idxprom997_3400_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom997_3400_resized;
      ov(13 downto 0) := iv;
      R_idxprom997_3400_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3401_index_1_resize
    process(idxprom997_3396) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom997_3396;
      ov := iv(13 downto 0);
      R_idxprom997_3400_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3401_root_address_inst
    process(array_obj_ref_3401_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3401_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3401_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3426_index_1_rename
    process(R_idxprom1002_3425_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1002_3425_resized;
      ov(13 downto 0) := iv;
      R_idxprom1002_3425_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3426_index_1_resize
    process(idxprom1002_3421) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1002_3421;
      ov := iv(13 downto 0);
      R_idxprom1002_3425_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3426_root_address_inst
    process(array_obj_ref_3426_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3426_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3426_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3898_index_1_rename
    process(R_idxprom1177_3897_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1177_3897_resized;
      ov(13 downto 0) := iv;
      R_idxprom1177_3897_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3898_index_1_resize
    process(idxprom1177_3893) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1177_3893;
      ov := iv(13 downto 0);
      R_idxprom1177_3897_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3898_root_address_inst
    process(array_obj_ref_3898_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3898_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3898_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3981_index_1_rename
    process(R_idxprom1220_3980_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1220_3980_resized;
      ov(13 downto 0) := iv;
      R_idxprom1220_3980_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3981_index_1_resize
    process(idxprom1220_3976) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1220_3976;
      ov := iv(13 downto 0);
      R_idxprom1220_3980_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3981_root_address_inst
    process(array_obj_ref_3981_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3981_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3981_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4006_index_1_rename
    process(R_idxprom1225_4005_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1225_4005_resized;
      ov(13 downto 0) := iv;
      R_idxprom1225_4005_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4006_index_1_resize
    process(idxprom1225_4001) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1225_4001;
      ov := iv(13 downto 0);
      R_idxprom1225_4005_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4006_root_address_inst
    process(array_obj_ref_4006_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4006_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4006_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4462_index_1_rename
    process(R_idxprom1395_4461_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1395_4461_resized;
      ov(13 downto 0) := iv;
      R_idxprom1395_4461_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4462_index_1_resize
    process(idxprom1395_4457) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1395_4457;
      ov := iv(13 downto 0);
      R_idxprom1395_4461_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4462_root_address_inst
    process(array_obj_ref_4462_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4462_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4462_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4545_index_1_rename
    process(R_idxprom1438_4544_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1438_4544_resized;
      ov(13 downto 0) := iv;
      R_idxprom1438_4544_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4545_index_1_resize
    process(idxprom1438_4540) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1438_4540;
      ov := iv(13 downto 0);
      R_idxprom1438_4544_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4545_root_address_inst
    process(array_obj_ref_4545_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4545_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4545_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4570_index_1_rename
    process(R_idxprom1443_4569_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1443_4569_resized;
      ov(13 downto 0) := iv;
      R_idxprom1443_4569_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4570_index_1_resize
    process(idxprom1443_4565) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1443_4565;
      ov := iv(13 downto 0);
      R_idxprom1443_4569_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_4570_root_address_inst
    process(array_obj_ref_4570_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_4570_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_4570_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5024_index_1_rename
    process(R_idxprom1615_5023_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1615_5023_resized;
      ov(13 downto 0) := iv;
      R_idxprom1615_5023_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5024_index_1_resize
    process(idxprom1615_5019) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1615_5019;
      ov := iv(13 downto 0);
      R_idxprom1615_5023_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5024_root_address_inst
    process(array_obj_ref_5024_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_5024_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_5024_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5107_index_1_rename
    process(R_idxprom1658_5106_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1658_5106_resized;
      ov(13 downto 0) := iv;
      R_idxprom1658_5106_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5107_index_1_resize
    process(idxprom1658_5102) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1658_5102;
      ov := iv(13 downto 0);
      R_idxprom1658_5106_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5107_root_address_inst
    process(array_obj_ref_5107_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_5107_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_5107_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5132_index_1_rename
    process(R_idxprom1663_5131_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1663_5131_resized;
      ov(13 downto 0) := iv;
      R_idxprom1663_5131_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5132_index_1_resize
    process(idxprom1663_5127) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1663_5127;
      ov := iv(13 downto 0);
      R_idxprom1663_5131_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_5132_root_address_inst
    process(array_obj_ref_5132_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_5132_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_5132_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_addr_0
    process(ptr_deref_1076_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1076_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_base_resize
    process(arrayidx_1074) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1074;
      ov := iv(13 downto 0);
      ptr_deref_1076_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_gather_scatter
    process(type_cast_1078_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1078_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1076_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1076_root_address_inst
    process(ptr_deref_1076_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1076_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1076_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_addr_0
    process(ptr_deref_1160_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1160_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_base_resize
    process(arrayidx131_1157) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx131_1157;
      ov := iv(13 downto 0);
      ptr_deref_1160_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_gather_scatter
    process(ptr_deref_1160_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_data_0;
      ov(63 downto 0) := iv;
      tmp132_1161 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1160_root_address_inst
    process(ptr_deref_1160_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1160_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1160_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_addr_0
    process(ptr_deref_1184_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1184_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1184_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_base_resize
    process(arrayidx136_1182) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx136_1182;
      ov := iv(13 downto 0);
      ptr_deref_1184_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_gather_scatter
    process(tmp132_1161) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp132_1161;
      ov(63 downto 0) := iv;
      ptr_deref_1184_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1184_root_address_inst
    process(ptr_deref_1184_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1184_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1184_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_addr_0
    process(ptr_deref_1359_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1359_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1359_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_base_resize
    process(iNsTr_22_1356) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_22_1356;
      ov := iv(6 downto 0);
      ptr_deref_1359_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_gather_scatter
    process(ptr_deref_1359_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1359_data_0;
      ov(31 downto 0) := iv;
      tmp213_1360 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_root_address_inst
    process(ptr_deref_1359_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1359_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1359_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_addr_0
    process(ptr_deref_1371_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1371_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1371_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_base_resize
    process(iNsTr_23_1368) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_23_1368;
      ov := iv(6 downto 0);
      ptr_deref_1371_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_gather_scatter
    process(ptr_deref_1371_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1371_data_0;
      ov(31 downto 0) := iv;
      tmp217_1372 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1371_root_address_inst
    process(ptr_deref_1371_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1371_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1371_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1632_addr_0
    process(ptr_deref_1632_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1632_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1632_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1632_base_resize
    process(arrayidx299_1630) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx299_1630;
      ov := iv(13 downto 0);
      ptr_deref_1632_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1632_gather_scatter
    process(type_cast_1634_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1634_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1632_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1632_root_address_inst
    process(ptr_deref_1632_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1632_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1632_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_addr_0
    process(ptr_deref_1716_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1716_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1716_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_base_resize
    process(arrayidx342_1713) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx342_1713;
      ov := iv(13 downto 0);
      ptr_deref_1716_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_gather_scatter
    process(ptr_deref_1716_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1716_data_0;
      ov(63 downto 0) := iv;
      tmp343_1717 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1716_root_address_inst
    process(ptr_deref_1716_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1716_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1716_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_addr_0
    process(ptr_deref_1740_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1740_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1740_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_base_resize
    process(arrayidx347_1738) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx347_1738;
      ov := iv(13 downto 0);
      ptr_deref_1740_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_gather_scatter
    process(tmp343_1717) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp343_1717;
      ov(63 downto 0) := iv;
      ptr_deref_1740_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1740_root_address_inst
    process(ptr_deref_1740_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1740_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1740_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_addr_0
    process(ptr_deref_1911_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1911_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1911_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_base_resize
    process(iNsTr_39_1908) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_1908;
      ov := iv(6 downto 0);
      ptr_deref_1911_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_gather_scatter
    process(ptr_deref_1911_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1911_data_0;
      ov(31 downto 0) := iv;
      tmp429_1912 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_root_address_inst
    process(ptr_deref_1911_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1911_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1911_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_addr_0
    process(ptr_deref_1923_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1923_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1923_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_base_resize
    process(iNsTr_40_1920) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_1920;
      ov := iv(6 downto 0);
      ptr_deref_1923_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_gather_scatter
    process(ptr_deref_1923_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1923_data_0;
      ov(31 downto 0) := iv;
      tmp433_1924 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_root_address_inst
    process(ptr_deref_1923_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1923_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1923_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2190_addr_0
    process(ptr_deref_2190_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2190_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2190_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2190_base_resize
    process(arrayidx516_2188) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx516_2188;
      ov := iv(13 downto 0);
      ptr_deref_2190_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2190_gather_scatter
    process(type_cast_2192_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2192_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2190_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2190_root_address_inst
    process(ptr_deref_2190_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2190_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2190_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2274_addr_0
    process(ptr_deref_2274_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2274_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2274_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2274_base_resize
    process(arrayidx559_2271) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx559_2271;
      ov := iv(13 downto 0);
      ptr_deref_2274_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2274_gather_scatter
    process(ptr_deref_2274_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2274_data_0;
      ov(63 downto 0) := iv;
      tmp560_2275 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2274_root_address_inst
    process(ptr_deref_2274_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2274_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2274_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_addr_0
    process(ptr_deref_2298_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2298_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2298_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_base_resize
    process(arrayidx564_2296) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx564_2296;
      ov := iv(13 downto 0);
      ptr_deref_2298_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_gather_scatter
    process(tmp560_2275) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp560_2275;
      ov(63 downto 0) := iv;
      ptr_deref_2298_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_root_address_inst
    process(ptr_deref_2298_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2298_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2298_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_addr_0
    process(ptr_deref_2486_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2486_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2486_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_base_resize
    process(iNsTr_56_2483) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_56_2483;
      ov := iv(6 downto 0);
      ptr_deref_2486_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_gather_scatter
    process(ptr_deref_2486_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2486_data_0;
      ov(31 downto 0) := iv;
      tmp651_2487 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_root_address_inst
    process(ptr_deref_2486_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2486_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2486_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_addr_0
    process(ptr_deref_2498_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2498_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2498_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_base_resize
    process(iNsTr_57_2495) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_57_2495;
      ov := iv(6 downto 0);
      ptr_deref_2498_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_gather_scatter
    process(ptr_deref_2498_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2498_data_0;
      ov(31 downto 0) := iv;
      tmp655_2499 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_root_address_inst
    process(ptr_deref_2498_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2498_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2498_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2758_addr_0
    process(ptr_deref_2758_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2758_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2758_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2758_base_resize
    process(arrayidx737_2756) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx737_2756;
      ov := iv(13 downto 0);
      ptr_deref_2758_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2758_gather_scatter
    process(type_cast_2760_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2760_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2758_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2758_root_address_inst
    process(ptr_deref_2758_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2758_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2758_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2842_addr_0
    process(ptr_deref_2842_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2842_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2842_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2842_base_resize
    process(arrayidx780_2839) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx780_2839;
      ov := iv(13 downto 0);
      ptr_deref_2842_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2842_gather_scatter
    process(ptr_deref_2842_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2842_data_0;
      ov(63 downto 0) := iv;
      tmp781_2843 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2842_root_address_inst
    process(ptr_deref_2842_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2842_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2842_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2866_addr_0
    process(ptr_deref_2866_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2866_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2866_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2866_base_resize
    process(arrayidx785_2864) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx785_2864;
      ov := iv(13 downto 0);
      ptr_deref_2866_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2866_gather_scatter
    process(tmp781_2843) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp781_2843;
      ov(63 downto 0) := iv;
      ptr_deref_2866_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2866_root_address_inst
    process(ptr_deref_2866_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2866_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2866_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3037_addr_0
    process(ptr_deref_3037_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3037_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3037_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3037_base_resize
    process(iNsTr_73_3034) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_73_3034;
      ov := iv(6 downto 0);
      ptr_deref_3037_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3037_gather_scatter
    process(ptr_deref_3037_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3037_data_0;
      ov(31 downto 0) := iv;
      tmp867_3038 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3037_root_address_inst
    process(ptr_deref_3037_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3037_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3037_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3049_addr_0
    process(ptr_deref_3049_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3049_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3049_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3049_base_resize
    process(iNsTr_74_3046) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_74_3046;
      ov := iv(6 downto 0);
      ptr_deref_3049_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3049_gather_scatter
    process(ptr_deref_3049_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3049_data_0;
      ov(31 downto 0) := iv;
      tmp871_3050 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3049_root_address_inst
    process(ptr_deref_3049_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3049_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3049_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3322_addr_0
    process(ptr_deref_3322_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3322_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3322_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3322_base_resize
    process(arrayidx955_3320) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx955_3320;
      ov := iv(13 downto 0);
      ptr_deref_3322_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3322_gather_scatter
    process(type_cast_3324_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3324_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3322_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3322_root_address_inst
    process(ptr_deref_3322_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3322_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3322_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3406_addr_0
    process(ptr_deref_3406_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3406_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3406_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3406_base_resize
    process(arrayidx998_3403) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx998_3403;
      ov := iv(13 downto 0);
      ptr_deref_3406_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3406_gather_scatter
    process(ptr_deref_3406_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3406_data_0;
      ov(63 downto 0) := iv;
      tmp999_3407 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3406_root_address_inst
    process(ptr_deref_3406_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3406_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3406_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3430_addr_0
    process(ptr_deref_3430_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3430_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3430_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3430_base_resize
    process(arrayidx1003_3428) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1003_3428;
      ov := iv(13 downto 0);
      ptr_deref_3430_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3430_gather_scatter
    process(tmp999_3407) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp999_3407;
      ov(63 downto 0) := iv;
      ptr_deref_3430_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3430_root_address_inst
    process(ptr_deref_3430_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3430_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3430_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3624_addr_0
    process(ptr_deref_3624_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3624_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3624_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3624_base_resize
    process(iNsTr_90_3621) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_90_3621;
      ov := iv(6 downto 0);
      ptr_deref_3624_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3624_gather_scatter
    process(ptr_deref_3624_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3624_data_0;
      ov(31 downto 0) := iv;
      tmp1091_3625 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3624_root_address_inst
    process(ptr_deref_3624_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3624_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3624_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_addr_0
    process(ptr_deref_3636_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3636_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_3636_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_base_resize
    process(iNsTr_91_3633) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_91_3633;
      ov := iv(6 downto 0);
      ptr_deref_3636_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_gather_scatter
    process(ptr_deref_3636_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3636_data_0;
      ov(31 downto 0) := iv;
      tmp1095_3637 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3636_root_address_inst
    process(ptr_deref_3636_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3636_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_3636_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3902_addr_0
    process(ptr_deref_3902_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3902_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3902_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3902_base_resize
    process(arrayidx1178_3900) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1178_3900;
      ov := iv(13 downto 0);
      ptr_deref_3902_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3902_gather_scatter
    process(type_cast_3904_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3904_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3902_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3902_root_address_inst
    process(ptr_deref_3902_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3902_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3902_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3986_addr_0
    process(ptr_deref_3986_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3986_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3986_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3986_base_resize
    process(arrayidx1221_3983) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1221_3983;
      ov := iv(13 downto 0);
      ptr_deref_3986_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3986_gather_scatter
    process(ptr_deref_3986_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3986_data_0;
      ov(63 downto 0) := iv;
      tmp1222_3987 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3986_root_address_inst
    process(ptr_deref_3986_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3986_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3986_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4010_addr_0
    process(ptr_deref_4010_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4010_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4010_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4010_base_resize
    process(arrayidx1226_4008) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1226_4008;
      ov := iv(13 downto 0);
      ptr_deref_4010_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4010_gather_scatter
    process(tmp1222_3987) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1222_3987;
      ov(63 downto 0) := iv;
      ptr_deref_4010_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4010_root_address_inst
    process(ptr_deref_4010_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4010_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4010_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4193_addr_0
    process(ptr_deref_4193_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4193_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4193_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4193_base_resize
    process(iNsTr_107_4190) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_107_4190;
      ov := iv(6 downto 0);
      ptr_deref_4193_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4193_gather_scatter
    process(ptr_deref_4193_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4193_data_0;
      ov(31 downto 0) := iv;
      tmp1310_4194 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4193_root_address_inst
    process(ptr_deref_4193_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4193_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4193_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_addr_0
    process(ptr_deref_4205_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4205_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4205_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_base_resize
    process(iNsTr_108_4202) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_108_4202;
      ov := iv(6 downto 0);
      ptr_deref_4205_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_gather_scatter
    process(ptr_deref_4205_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4205_data_0;
      ov(31 downto 0) := iv;
      tmp1314_4206 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4205_root_address_inst
    process(ptr_deref_4205_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4205_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4205_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4466_addr_0
    process(ptr_deref_4466_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4466_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4466_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4466_base_resize
    process(arrayidx1396_4464) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1396_4464;
      ov := iv(13 downto 0);
      ptr_deref_4466_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4466_gather_scatter
    process(type_cast_4468_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_4468_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_4466_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4466_root_address_inst
    process(ptr_deref_4466_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4466_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4466_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4550_addr_0
    process(ptr_deref_4550_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4550_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4550_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4550_base_resize
    process(arrayidx1439_4547) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1439_4547;
      ov := iv(13 downto 0);
      ptr_deref_4550_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4550_gather_scatter
    process(ptr_deref_4550_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4550_data_0;
      ov(63 downto 0) := iv;
      tmp1440_4551 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4550_root_address_inst
    process(ptr_deref_4550_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4550_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4550_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4574_addr_0
    process(ptr_deref_4574_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4574_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_4574_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4574_base_resize
    process(arrayidx1444_4572) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1444_4572;
      ov := iv(13 downto 0);
      ptr_deref_4574_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4574_gather_scatter
    process(tmp1440_4551) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1440_4551;
      ov(63 downto 0) := iv;
      ptr_deref_4574_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4574_root_address_inst
    process(ptr_deref_4574_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4574_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_4574_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4762_addr_0
    process(ptr_deref_4762_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4762_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4762_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4762_base_resize
    process(iNsTr_124_4759) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_124_4759;
      ov := iv(6 downto 0);
      ptr_deref_4762_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4762_gather_scatter
    process(ptr_deref_4762_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4762_data_0;
      ov(31 downto 0) := iv;
      tmp1531_4763 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4762_root_address_inst
    process(ptr_deref_4762_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4762_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4762_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4774_addr_0
    process(ptr_deref_4774_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4774_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_4774_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4774_base_resize
    process(iNsTr_125_4771) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_125_4771;
      ov := iv(6 downto 0);
      ptr_deref_4774_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4774_gather_scatter
    process(ptr_deref_4774_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4774_data_0;
      ov(31 downto 0) := iv;
      tmp1535_4775 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_4774_root_address_inst
    process(ptr_deref_4774_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_4774_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_4774_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5028_addr_0
    process(ptr_deref_5028_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5028_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_5028_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5028_base_resize
    process(arrayidx1616_5026) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1616_5026;
      ov := iv(13 downto 0);
      ptr_deref_5028_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5028_gather_scatter
    process(type_cast_5030_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_5030_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_5028_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5028_root_address_inst
    process(ptr_deref_5028_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5028_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_5028_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5112_addr_0
    process(ptr_deref_5112_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5112_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_5112_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5112_base_resize
    process(arrayidx1659_5109) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1659_5109;
      ov := iv(13 downto 0);
      ptr_deref_5112_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5112_gather_scatter
    process(ptr_deref_5112_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5112_data_0;
      ov(63 downto 0) := iv;
      tmp1660_5113 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5112_root_address_inst
    process(ptr_deref_5112_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5112_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_5112_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5136_addr_0
    process(ptr_deref_5136_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5136_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_5136_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5136_base_resize
    process(arrayidx1664_5134) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1664_5134;
      ov := iv(13 downto 0);
      ptr_deref_5136_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5136_gather_scatter
    process(tmp1660_5113) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1660_5113;
      ov(63 downto 0) := iv;
      ptr_deref_5136_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_5136_root_address_inst
    process(ptr_deref_5136_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_5136_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_5136_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_addr_0
    process(ptr_deref_727_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_727_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_base_resize
    process(iNsTr_0_724) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_724;
      ov := iv(6 downto 0);
      ptr_deref_727_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_gather_scatter
    process(ptr_deref_727_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_data_0;
      ov(31 downto 0) := iv;
      tmp_728 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_727_root_address_inst
    process(ptr_deref_727_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_727_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_727_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_addr_0
    process(ptr_deref_746_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_746_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_746_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_base_resize
    process(iNsTr_2_743) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_743;
      ov := iv(6 downto 0);
      ptr_deref_746_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_gather_scatter
    process(ptr_deref_746_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_746_data_0;
      ov(31 downto 0) := iv;
      tmp1_747 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_746_root_address_inst
    process(ptr_deref_746_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_746_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_746_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_addr_0
    process(ptr_deref_765_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_765_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_765_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_base_resize
    process(iNsTr_4_762) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_762;
      ov := iv(6 downto 0);
      ptr_deref_765_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_gather_scatter
    process(ptr_deref_765_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_765_data_0;
      ov(31 downto 0) := iv;
      tmp3_766 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_765_root_address_inst
    process(ptr_deref_765_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_765_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_765_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_addr_0
    process(ptr_deref_794_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_794_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_794_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_base_resize
    process(iNsTr_7_791) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_791;
      ov := iv(6 downto 0);
      ptr_deref_794_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_gather_scatter
    process(ptr_deref_794_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_794_data_0;
      ov(31 downto 0) := iv;
      tmp21_795 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_794_root_address_inst
    process(ptr_deref_794_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_794_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_794_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_addr_0
    process(ptr_deref_806_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_806_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_806_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_base_resize
    process(iNsTr_8_803) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_803;
      ov := iv(6 downto 0);
      ptr_deref_806_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_gather_scatter
    process(ptr_deref_806_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_806_data_0;
      ov(31 downto 0) := iv;
      tmp24_807 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_806_root_address_inst
    process(ptr_deref_806_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_806_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_806_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1016_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp74_1015;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1016_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1016_branch_req_0,
          ack0 => if_stmt_1016_branch_ack_0,
          ack1 => if_stmt_1016_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1207_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp143_1206;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1207_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1207_branch_req_0,
          ack0 => if_stmt_1207_branch_ack_0,
          ack1 => if_stmt_1207_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1300_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp176_1299;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1300_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1300_branch_req_0,
          ack0 => if_stmt_1300_branch_ack_0,
          ack1 => if_stmt_1300_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1496_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp249_1495;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1496_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1496_branch_req_0,
          ack0 => if_stmt_1496_branch_ack_0,
          ack1 => if_stmt_1496_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1528_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp260_1527;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1528_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1528_branch_req_0,
          ack0 => if_stmt_1528_branch_ack_0,
          ack1 => if_stmt_1528_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1547_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp267_1546;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1547_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1547_branch_req_0,
          ack0 => if_stmt_1547_branch_ack_0,
          ack1 => if_stmt_1547_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1573_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp277_1572;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1573_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1573_branch_req_0,
          ack0 => if_stmt_1573_branch_ack_0,
          ack1 => if_stmt_1573_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1763_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp356_1762;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1763_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1763_branch_req_0,
          ack0 => if_stmt_1763_branch_ack_0,
          ack1 => if_stmt_1763_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1849_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp390_1848;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1849_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1849_branch_req_0,
          ack0 => if_stmt_1849_branch_ack_0,
          ack1 => if_stmt_1849_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2048_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp465_2047;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2048_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2048_branch_req_0,
          ack0 => if_stmt_2048_branch_ack_0,
          ack1 => if_stmt_2048_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2080_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp476_2079;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2080_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2080_branch_req_0,
          ack0 => if_stmt_2080_branch_ack_0,
          ack1 => if_stmt_2080_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2099_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp483_2098;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2099_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2099_branch_req_0,
          ack0 => if_stmt_2099_branch_ack_0,
          ack1 => if_stmt_2099_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2131_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp494_2130;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2131_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2131_branch_req_0,
          ack0 => if_stmt_2131_branch_ack_0,
          ack1 => if_stmt_2131_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2321_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp573_2320;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2321_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2321_branch_req_0,
          ack0 => if_stmt_2321_branch_ack_0,
          ack1 => if_stmt_2321_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2414_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp608_2413;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2414_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2414_branch_req_0,
          ack0 => if_stmt_2414_branch_ack_0,
          ack1 => if_stmt_2414_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2622_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp687_2621;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2622_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2622_branch_req_0,
          ack0 => if_stmt_2622_branch_ack_0,
          ack1 => if_stmt_2622_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2654_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp698_2653;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2654_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2654_branch_req_0,
          ack0 => if_stmt_2654_branch_ack_0,
          ack1 => if_stmt_2654_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2673_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp705_2672;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2673_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2673_branch_req_0,
          ack0 => if_stmt_2673_branch_ack_0,
          ack1 => if_stmt_2673_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2699_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp715_2698;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2699_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2699_branch_req_0,
          ack0 => if_stmt_2699_branch_ack_0,
          ack1 => if_stmt_2699_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2889_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp794_2888;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2889_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2889_branch_req_0,
          ack0 => if_stmt_2889_branch_ack_0,
          ack1 => if_stmt_2889_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2975_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp828_2974;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2975_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2975_branch_req_0,
          ack0 => if_stmt_2975_branch_ack_0,
          ack1 => if_stmt_2975_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3174_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp903_3173;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3174_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3174_branch_req_0,
          ack0 => if_stmt_3174_branch_ack_0,
          ack1 => if_stmt_3174_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3212_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp915_3211;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3212_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3212_branch_req_0,
          ack0 => if_stmt_3212_branch_ack_0,
          ack1 => if_stmt_3212_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3231_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp922_3230;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3231_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3231_branch_req_0,
          ack0 => if_stmt_3231_branch_ack_0,
          ack1 => if_stmt_3231_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3263_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp933_3262;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3263_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3263_branch_req_0,
          ack0 => if_stmt_3263_branch_ack_0,
          ack1 => if_stmt_3263_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3453_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1012_3452;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3453_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3453_branch_req_0,
          ack0 => if_stmt_3453_branch_ack_0,
          ack1 => if_stmt_3453_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3552_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1048_3551;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3552_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3552_branch_req_0,
          ack0 => if_stmt_3552_branch_ack_0,
          ack1 => if_stmt_3552_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3760_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1127_3759;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3760_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3760_branch_req_0,
          ack0 => if_stmt_3760_branch_ack_0,
          ack1 => if_stmt_3760_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3798_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1139_3797;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3798_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3798_branch_req_0,
          ack0 => if_stmt_3798_branch_ack_0,
          ack1 => if_stmt_3798_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3817_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1146_3816;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3817_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3817_branch_req_0,
          ack0 => if_stmt_3817_branch_ack_0,
          ack1 => if_stmt_3817_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3843_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1156_3842;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3843_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3843_branch_req_0,
          ack0 => if_stmt_3843_branch_ack_0,
          ack1 => if_stmt_3843_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4033_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1235_4032;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4033_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4033_branch_req_0,
          ack0 => if_stmt_4033_branch_ack_0,
          ack1 => if_stmt_4033_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4125_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1270_4124;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4125_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4125_branch_req_0,
          ack0 => if_stmt_4125_branch_ack_0,
          ack1 => if_stmt_4125_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4330_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1346_4329;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4330_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4330_branch_req_0,
          ack0 => if_stmt_4330_branch_ack_0,
          ack1 => if_stmt_4330_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4356_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1356_4355;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4356_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4356_branch_req_0,
          ack0 => if_stmt_4356_branch_ack_0,
          ack1 => if_stmt_4356_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4375_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1363_4374;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4375_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4375_branch_req_0,
          ack0 => if_stmt_4375_branch_ack_0,
          ack1 => if_stmt_4375_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4407_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1374_4406;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4407_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4407_branch_req_0,
          ack0 => if_stmt_4407_branch_ack_0,
          ack1 => if_stmt_4407_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4597_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1453_4596;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4597_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4597_branch_req_0,
          ack0 => if_stmt_4597_branch_ack_0,
          ack1 => if_stmt_4597_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4684_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1487_4683;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4684_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4684_branch_req_0,
          ack0 => if_stmt_4684_branch_ack_0,
          ack1 => if_stmt_4684_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4898_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1567_4897;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4898_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4898_branch_req_0,
          ack0 => if_stmt_4898_branch_ack_0,
          ack1 => if_stmt_4898_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4924_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1577_4923;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4924_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4924_branch_req_0,
          ack0 => if_stmt_4924_branch_ack_0,
          ack1 => if_stmt_4924_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4943_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1584_4942;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4943_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4943_branch_req_0,
          ack0 => if_stmt_4943_branch_ack_0,
          ack1 => if_stmt_4943_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_4969_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1594_4968;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_4969_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_4969_branch_req_0,
          ack0 => if_stmt_4969_branch_ack_0,
          ack1 => if_stmt_4969_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_5159_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1673_5158;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_5159_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_5159_branch_req_0,
          ack0 => if_stmt_5159_branch_ack_0,
          ack1 => if_stmt_5159_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_5239_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1706_5238;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_5239_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_5239_branch_req_0,
          ack0 => if_stmt_5239_branch_ack_0,
          ack1 => if_stmt_5239_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_933_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_932;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_933_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_933_branch_req_0,
          ack0 => if_stmt_933_branch_ack_0,
          ack1 => if_stmt_933_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_965_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp56_964;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_965_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_965_branch_req_0,
          ack0 => if_stmt_965_branch_ack_0,
          ack1 => if_stmt_965_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_984_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp63_983;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_984_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_984_branch_req_0,
          ack0 => if_stmt_984_branch_ack_0,
          ack1 => if_stmt_984_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1218_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_913, type_cast_1217_wire_constant, tmp_var);
      add148_1219 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1226_inst
    process(jx_x1_899) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_899, type_cast_1225_wire_constant, tmp_var);
      inc_1227 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1263_inst
    process(inc165_1259, ix_x2_906) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc165_1259, ix_x2_906, tmp_var);
      inc165x_xix_x2_1264 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1774_inst
    process(k186x_x1_1476) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k186x_x1_1476, type_cast_1773_wire_constant, tmp_var);
      add361_1775 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1782_inst
    process(j240x_x1_1463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j240x_x1_1463, type_cast_1781_wire_constant, tmp_var);
      inc365_1783 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1813_inst
    process(inc379_1809, i194x_x2_1469) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc379_1809, i194x_x2_1469, tmp_var);
      inc379x_xi194x_x2_1814 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2332_inst
    process(k402x_x1_2015) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k402x_x1_2015, type_cast_2331_wire_constant, tmp_var);
      add578_2333 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2340_inst
    process(j456x_x1_2028) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j456x_x1_2028, type_cast_2339_wire_constant, tmp_var);
      inc582_2341 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2377_inst
    process(inc597_2373, i406x_x2_2022) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc597_2373, i406x_x2_2022, tmp_var);
      inc597x_xi406x_x2_2378 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2900_inst
    process(k620x_x1_2590) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k620x_x1_2590, type_cast_2899_wire_constant, tmp_var);
      add799_2901 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2908_inst
    process(j678x_x1_2603) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j678x_x1_2603, type_cast_2907_wire_constant, tmp_var);
      inc803_2909 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2939_inst
    process(inc817_2935, i628x_x2_2597) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc817_2935, i628x_x2_2597, tmp_var);
      inc817x_xi628x_x2_2940 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3464_inst
    process(k840x_x1_3141) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k840x_x1_3141, type_cast_3463_wire_constant, tmp_var);
      add1017_3465 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3472_inst
    process(j894x_x1_3154) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j894x_x1_3154, type_cast_3471_wire_constant, tmp_var);
      inc1021_3473 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3509_inst
    process(inc1036_3505, i844x_x2_3148) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1036_3505, i844x_x2_3148, tmp_var);
      inc1036x_xi844x_x2_3510 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4044_inst
    process(k1060x_x1_3728) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1060x_x1_3728, type_cast_4043_wire_constant, tmp_var);
      add1240_4045 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4052_inst
    process(j1118x_x1_3741) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1118x_x1_3741, type_cast_4051_wire_constant, tmp_var);
      inc1244_4053 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4083_inst
    process(inc1258_4079, i1068x_x2_3735) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1258_4079, i1068x_x2_3735, tmp_var);
      inc1258x_xi1068x_x2_4084 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4608_inst
    process(k1282x_x1_4297) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1282x_x1_4297, type_cast_4607_wire_constant, tmp_var);
      add1458_4609 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4616_inst
    process(j1337x_x1_4310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1337x_x1_4310, type_cast_4615_wire_constant, tmp_var);
      inc1462_4617 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_4653_inst
    process(inc1477_4649, i1286x_x2_4304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1477_4649, i1286x_x2_4304, tmp_var);
      inc1477x_xi1286x_x2_4654 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_5170_inst
    process(k1499x_x1_4866) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1499x_x1_4866, type_cast_5169_wire_constant, tmp_var);
      add1678_5171 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_5178_inst
    process(j1558x_x1_4879) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1558x_x1_4879, type_cast_5177_wire_constant, tmp_var);
      inc1682_5179 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_5209_inst
    process(inc1696_5205, i1507x_x2_4873) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1696_5205, i1507x_x2_4873, tmp_var);
      inc1696x_xi1507x_x2_5210 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1007_inst
    process(div70_1003, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div70_1003, conv48_855, tmp_var);
      add73_1008 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1046_inst
    process(mul89_1042, mul83_1037) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul89_1042, mul83_1037, tmp_var);
      add84_1047 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1051_inst
    process(add84_1047, conv78_1027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add84_1047, conv78_1027, tmp_var);
      add90_1052 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1110_inst
    process(conv94_1086, mul101_1096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv94_1086, mul101_1096, tmp_var);
      add102_1111 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1115_inst
    process(add102_1111, mul110_1106) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add102_1111, mul110_1106, tmp_var);
      add111_1116 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1130_inst
    process(mul126_1126, mul120_1121) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul126_1126, mul120_1121, tmp_var);
      add121_1131 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1135_inst
    process(add121_1131, conv94_1086) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add121_1131, conv94_1086, tmp_var);
      add127_1136 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1198_inst
    process(conv139_1193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv139_1193, type_cast_1197_wire_constant, tmp_var);
      add140_1199 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1249_inst
    process(div156_1245, shl_876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div156_1245, shl_876, tmp_var);
      add159_1250 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1293_inst
    process(div171_1289, shl_876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div171_1289, shl_876, tmp_var);
      add175_1294 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1519_inst
    process(div256_1515, conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div256_1515, conv248_1419, tmp_var);
      add259_1520 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1564_inst
    process(conv273_1560, conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv273_1560, conv248_1419, tmp_var);
      add276_1565 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1603_inst
    process(mul294_1599, mul288_1594) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul294_1599, mul288_1594, tmp_var);
      add289_1604 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1608_inst
    process(add289_1604, conv283_1584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add289_1604, conv283_1584, tmp_var);
      add295_1609 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1666_inst
    process(conv304_1642, mul312_1652) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv304_1642, mul312_1652, tmp_var);
      add313_1667 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1671_inst
    process(add313_1667, mul321_1662) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add313_1667, mul321_1662, tmp_var);
      add322_1672 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1686_inst
    process(mul337_1682, mul331_1677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul337_1682, mul331_1677, tmp_var);
      add332_1687 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1691_inst
    process(add332_1687, conv304_1642) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add332_1687, conv304_1642, tmp_var);
      add338_1692 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1754_inst
    process(conv352_1749) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv352_1749, type_cast_1753_wire_constant, tmp_var);
      add353_1755 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1799_inst
    process(conv369_1795, shl372_1440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv369_1795, shl372_1440, tmp_var);
      add373_1800 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1842_inst
    process(div385_1838, shl372_1440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div385_1838, shl372_1440, tmp_var);
      add389_1843 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2071_inst
    process(div472_2067, conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div472_2067, conv464_1971, tmp_var);
      add475_2072 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2122_inst
    process(div490_2118, conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div490_2118, conv464_1971, tmp_var);
      add493_2123 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2161_inst
    process(mul511_2157, conv500_2142) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul511_2157, conv500_2142, tmp_var);
      add506_2162 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2166_inst
    process(add506_2162, mul505_2152) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add506_2162, mul505_2152, tmp_var);
      add512_2167 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2224_inst
    process(mul538_2220, conv521_2200) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul538_2220, conv521_2200, tmp_var);
      add530_2225 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2229_inst
    process(add530_2225, mul529_2210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add530_2225, mul529_2210, tmp_var);
      add539_2230 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2244_inst
    process(mul554_2240, conv521_2200) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul554_2240, conv521_2200, tmp_var);
      add549_2245 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2249_inst
    process(add549_2245, mul548_2235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add549_2245, mul548_2235, tmp_var);
      add555_2250 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2312_inst
    process(conv569_2307) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv569_2307, type_cast_2311_wire_constant, tmp_var);
      add570_2313 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2363_inst
    process(div587_2359, shl590_1992) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div587_2359, shl590_1992, tmp_var);
      add591_2364 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2407_inst
    process(div603_2403, shl590_1992) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div603_2403, shl590_1992, tmp_var);
      add607_2408 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2645_inst
    process(div694_2641, conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div694_2641, conv686_2546, tmp_var);
      add697_2646 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2690_inst
    process(conv711_2686, conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv711_2686, conv686_2546, tmp_var);
      add714_2691 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2729_inst
    process(mul732_2725, conv721_2710) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul732_2725, conv721_2710, tmp_var);
      add727_2730 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2734_inst
    process(add727_2730, mul726_2720) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add727_2730, mul726_2720, tmp_var);
      add733_2735 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2792_inst
    process(mul759_2788, conv742_2768) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul759_2788, conv742_2768, tmp_var);
      add751_2793 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2797_inst
    process(add751_2793, mul750_2778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add751_2793, mul750_2778, tmp_var);
      add760_2798 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2812_inst
    process(mul775_2808, conv742_2768) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul775_2808, conv742_2768, tmp_var);
      add770_2813 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2817_inst
    process(add770_2813, mul769_2803) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add770_2813, mul769_2803, tmp_var);
      add776_2818 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2880_inst
    process(conv790_2875) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv790_2875, type_cast_2879_wire_constant, tmp_var);
      add791_2881 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2925_inst
    process(conv807_2921, shl810_2567) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv807_2921, shl810_2567, tmp_var);
      add811_2926 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2968_inst
    process(div823_2964, shl810_2567) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div823_2964, shl810_2567, tmp_var);
      add827_2969 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3203_inst
    process(div911_3199, conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div911_3199, conv902_3097, tmp_var);
      add914_3204 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3254_inst
    process(div929_3250, conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div929_3250, conv902_3097, tmp_var);
      add932_3255 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3293_inst
    process(mul950_3289, conv939_3274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul950_3289, conv939_3274, tmp_var);
      add945_3294 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3298_inst
    process(add945_3294, mul944_3284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add945_3294, mul944_3284, tmp_var);
      add951_3299 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3356_inst
    process(mul977_3352, conv960_3332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul977_3352, conv960_3332, tmp_var);
      add969_3357 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3361_inst
    process(add969_3357, mul968_3342) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add969_3357, mul968_3342, tmp_var);
      add978_3362 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3376_inst
    process(mul993_3372, conv960_3332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul993_3372, conv960_3332, tmp_var);
      add988_3377 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3381_inst
    process(add988_3377, mul987_3367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add988_3377, mul987_3367, tmp_var);
      add994_3382 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3444_inst
    process(conv1008_3439) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1008_3439, type_cast_3443_wire_constant, tmp_var);
      add1009_3445 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3495_inst
    process(div1026_3491, shl1029_3118) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1026_3491, shl1029_3118, tmp_var);
      add1030_3496 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3545_inst
    process(div1043_3541, shl1029_3118) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1043_3541, shl1029_3118, tmp_var);
      add1047_3546 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3789_inst
    process(div1135_3785, conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1135_3785, conv1126_3684, tmp_var);
      add1138_3790 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3834_inst
    process(conv1152_3830, conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1152_3830, conv1126_3684, tmp_var);
      add1155_3835 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3873_inst
    process(mul1173_3869, conv1162_3854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1173_3869, conv1162_3854, tmp_var);
      add1168_3874 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3878_inst
    process(add1168_3874, mul1167_3864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1168_3874, mul1167_3864, tmp_var);
      add1174_3879 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3936_inst
    process(mul1200_3932, conv1183_3912) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1200_3932, conv1183_3912, tmp_var);
      add1192_3937 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3941_inst
    process(add1192_3937, mul1191_3922) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1192_3937, mul1191_3922, tmp_var);
      add1201_3942 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3956_inst
    process(mul1216_3952, conv1183_3912) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1216_3952, conv1183_3912, tmp_var);
      add1211_3957 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3961_inst
    process(add1211_3957, mul1210_3947) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1211_3957, mul1210_3947, tmp_var);
      add1217_3962 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4024_inst
    process(conv1231_4019) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1231_4019, type_cast_4023_wire_constant, tmp_var);
      add1232_4025 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4069_inst
    process(conv1248_4065, shl1251_3705) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1248_4065, shl1251_3705, tmp_var);
      add1252_4070 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4118_inst
    process(div1265_4114, shl1251_3705) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1265_4114, shl1251_3705, tmp_var);
      add1269_4119 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4347_inst
    process(conv1352_4343, conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1352_4343, conv1345_4253, tmp_var);
      add1355_4348 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4398_inst
    process(div1370_4394, conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1370_4394, conv1345_4253, tmp_var);
      add1373_4399 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4437_inst
    process(mul1391_4433, conv1380_4418) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1391_4433, conv1380_4418, tmp_var);
      add1386_4438 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4442_inst
    process(add1386_4438, mul1385_4428) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1386_4438, mul1385_4428, tmp_var);
      add1392_4443 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4500_inst
    process(mul1418_4496, conv1401_4476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1418_4496, conv1401_4476, tmp_var);
      add1410_4501 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4505_inst
    process(add1410_4501, mul1409_4486) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1410_4501, mul1409_4486, tmp_var);
      add1419_4506 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4520_inst
    process(mul1434_4516, conv1401_4476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1434_4516, conv1401_4476, tmp_var);
      add1429_4521 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4525_inst
    process(add1429_4521, mul1428_4511) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1429_4521, mul1428_4511, tmp_var);
      add1435_4526 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4588_inst
    process(conv1449_4583) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1449_4583, type_cast_4587_wire_constant, tmp_var);
      add1450_4589 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4639_inst
    process(div1467_4635, shl1470_4274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div1467_4635, shl1470_4274, tmp_var);
      add1471_4640 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4677_inst
    process(conv1482_4673, shl1470_4274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1482_4673, shl1470_4274, tmp_var);
      add1486_4678 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4915_inst
    process(conv1573_4911, conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1573_4911, conv1566_4822, tmp_var);
      add1576_4916 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4960_inst
    process(conv1590_4956, conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1590_4956, conv1566_4822, tmp_var);
      add1593_4961 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_4999_inst
    process(mul1611_4995, conv1600_4980) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1611_4995, conv1600_4980, tmp_var);
      add1606_5000 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5004_inst
    process(add1606_5000, mul1605_4990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1606_5000, mul1605_4990, tmp_var);
      add1612_5005 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5062_inst
    process(mul1638_5058, conv1621_5038) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1638_5058, conv1621_5038, tmp_var);
      add1630_5063 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5067_inst
    process(add1630_5063, mul1629_5048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1630_5063, mul1629_5048, tmp_var);
      add1639_5068 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5082_inst
    process(mul1654_5078, conv1621_5038) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1654_5078, conv1621_5038, tmp_var);
      add1649_5083 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5087_inst
    process(add1649_5083, mul1648_5073) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1649_5083, mul1648_5073, tmp_var);
      add1655_5088 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5150_inst
    process(conv1669_5145) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1669_5145, type_cast_5149_wire_constant, tmp_var);
      add1670_5151 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5195_inst
    process(conv1686_5191, shl1689_4843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1686_5191, shl1689_4843, tmp_var);
      add1690_5196 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_5232_inst
    process(conv1701_5228, shl1689_4843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1701_5228, shl1689_4843, tmp_var);
      add1705_5233 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_956_inst
    process(div_952, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(div_952, conv48_855, tmp_var);
      add_957 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1059_inst
    process(type_cast_1055_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1055_wire, type_cast_1058_wire_constant, tmp_var);
      ASHR_i32_i32_1059_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1143_inst
    process(type_cast_1139_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1139_wire, type_cast_1142_wire_constant, tmp_var);
      ASHR_i32_i32_1143_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1168_inst
    process(type_cast_1164_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1164_wire, type_cast_1167_wire_constant, tmp_var);
      ASHR_i32_i32_1168_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1393_inst
    process(type_cast_1389_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1389_wire, type_cast_1392_wire_constant, tmp_var);
      ASHR_i32_i32_1393_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1408_inst
    process(type_cast_1404_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1404_wire, type_cast_1407_wire_constant, tmp_var);
      ASHR_i32_i32_1408_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1432_inst
    process(type_cast_1428_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1428_wire, type_cast_1431_wire_constant, tmp_var);
      ASHR_i32_i32_1432_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1458_inst
    process(type_cast_1454_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1454_wire, type_cast_1457_wire_constant, tmp_var);
      ASHR_i32_i32_1458_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1616_inst
    process(type_cast_1612_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1612_wire, type_cast_1615_wire_constant, tmp_var);
      ASHR_i32_i32_1616_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1699_inst
    process(type_cast_1695_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1695_wire, type_cast_1698_wire_constant, tmp_var);
      ASHR_i32_i32_1699_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1724_inst
    process(type_cast_1720_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1720_wire, type_cast_1723_wire_constant, tmp_var);
      ASHR_i32_i32_1724_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1945_inst
    process(type_cast_1941_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1941_wire, type_cast_1944_wire_constant, tmp_var);
      ASHR_i32_i32_1945_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1960_inst
    process(type_cast_1956_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1956_wire, type_cast_1959_wire_constant, tmp_var);
      ASHR_i32_i32_1960_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1984_inst
    process(type_cast_1980_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1980_wire, type_cast_1983_wire_constant, tmp_var);
      ASHR_i32_i32_1984_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2010_inst
    process(type_cast_2006_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2006_wire, type_cast_2009_wire_constant, tmp_var);
      ASHR_i32_i32_2010_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2174_inst
    process(type_cast_2170_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2170_wire, type_cast_2173_wire_constant, tmp_var);
      ASHR_i32_i32_2174_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2257_inst
    process(type_cast_2253_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2253_wire, type_cast_2256_wire_constant, tmp_var);
      ASHR_i32_i32_2257_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2282_inst
    process(type_cast_2278_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2278_wire, type_cast_2281_wire_constant, tmp_var);
      ASHR_i32_i32_2282_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2520_inst
    process(type_cast_2516_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2516_wire, type_cast_2519_wire_constant, tmp_var);
      ASHR_i32_i32_2520_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2535_inst
    process(type_cast_2531_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2531_wire, type_cast_2534_wire_constant, tmp_var);
      ASHR_i32_i32_2535_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2559_inst
    process(type_cast_2555_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2555_wire, type_cast_2558_wire_constant, tmp_var);
      ASHR_i32_i32_2559_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2585_inst
    process(type_cast_2581_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2581_wire, type_cast_2584_wire_constant, tmp_var);
      ASHR_i32_i32_2585_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2742_inst
    process(type_cast_2738_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2738_wire, type_cast_2741_wire_constant, tmp_var);
      ASHR_i32_i32_2742_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2825_inst
    process(type_cast_2821_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2821_wire, type_cast_2824_wire_constant, tmp_var);
      ASHR_i32_i32_2825_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2850_inst
    process(type_cast_2846_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2846_wire, type_cast_2849_wire_constant, tmp_var);
      ASHR_i32_i32_2850_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3071_inst
    process(type_cast_3067_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3067_wire, type_cast_3070_wire_constant, tmp_var);
      ASHR_i32_i32_3071_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3086_inst
    process(type_cast_3082_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3082_wire, type_cast_3085_wire_constant, tmp_var);
      ASHR_i32_i32_3086_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3110_inst
    process(type_cast_3106_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3106_wire, type_cast_3109_wire_constant, tmp_var);
      ASHR_i32_i32_3110_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3136_inst
    process(type_cast_3132_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3132_wire, type_cast_3135_wire_constant, tmp_var);
      ASHR_i32_i32_3136_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3306_inst
    process(type_cast_3302_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3302_wire, type_cast_3305_wire_constant, tmp_var);
      ASHR_i32_i32_3306_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3389_inst
    process(type_cast_3385_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3385_wire, type_cast_3388_wire_constant, tmp_var);
      ASHR_i32_i32_3389_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3414_inst
    process(type_cast_3410_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3410_wire, type_cast_3413_wire_constant, tmp_var);
      ASHR_i32_i32_3414_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3658_inst
    process(type_cast_3654_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3654_wire, type_cast_3657_wire_constant, tmp_var);
      ASHR_i32_i32_3658_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3673_inst
    process(type_cast_3669_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3669_wire, type_cast_3672_wire_constant, tmp_var);
      ASHR_i32_i32_3673_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3697_inst
    process(type_cast_3693_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3693_wire, type_cast_3696_wire_constant, tmp_var);
      ASHR_i32_i32_3697_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3723_inst
    process(type_cast_3719_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3719_wire, type_cast_3722_wire_constant, tmp_var);
      ASHR_i32_i32_3723_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3886_inst
    process(type_cast_3882_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3882_wire, type_cast_3885_wire_constant, tmp_var);
      ASHR_i32_i32_3886_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3969_inst
    process(type_cast_3965_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3965_wire, type_cast_3968_wire_constant, tmp_var);
      ASHR_i32_i32_3969_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3994_inst
    process(type_cast_3990_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3990_wire, type_cast_3993_wire_constant, tmp_var);
      ASHR_i32_i32_3994_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4227_inst
    process(type_cast_4223_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4223_wire, type_cast_4226_wire_constant, tmp_var);
      ASHR_i32_i32_4227_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4242_inst
    process(type_cast_4238_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4238_wire, type_cast_4241_wire_constant, tmp_var);
      ASHR_i32_i32_4242_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4266_inst
    process(type_cast_4262_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4262_wire, type_cast_4265_wire_constant, tmp_var);
      ASHR_i32_i32_4266_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4292_inst
    process(type_cast_4288_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4288_wire, type_cast_4291_wire_constant, tmp_var);
      ASHR_i32_i32_4292_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4450_inst
    process(type_cast_4446_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4446_wire, type_cast_4449_wire_constant, tmp_var);
      ASHR_i32_i32_4450_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4533_inst
    process(type_cast_4529_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4529_wire, type_cast_4532_wire_constant, tmp_var);
      ASHR_i32_i32_4533_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4558_inst
    process(type_cast_4554_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4554_wire, type_cast_4557_wire_constant, tmp_var);
      ASHR_i32_i32_4558_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4796_inst
    process(type_cast_4792_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4792_wire, type_cast_4795_wire_constant, tmp_var);
      ASHR_i32_i32_4796_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4811_inst
    process(type_cast_4807_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4807_wire, type_cast_4810_wire_constant, tmp_var);
      ASHR_i32_i32_4811_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4835_inst
    process(type_cast_4831_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4831_wire, type_cast_4834_wire_constant, tmp_var);
      ASHR_i32_i32_4835_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_4861_inst
    process(type_cast_4857_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_4857_wire, type_cast_4860_wire_constant, tmp_var);
      ASHR_i32_i32_4861_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_5012_inst
    process(type_cast_5008_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_5008_wire, type_cast_5011_wire_constant, tmp_var);
      ASHR_i32_i32_5012_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_5095_inst
    process(type_cast_5091_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_5091_wire, type_cast_5094_wire_constant, tmp_var);
      ASHR_i32_i32_5095_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_5120_inst
    process(type_cast_5116_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_5116_wire, type_cast_5119_wire_constant, tmp_var);
      ASHR_i32_i32_5120_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_829_inst
    process(type_cast_825_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_825_wire, type_cast_828_wire_constant, tmp_var);
      ASHR_i32_i32_829_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_844_inst
    process(type_cast_840_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_840_wire, type_cast_843_wire_constant, tmp_var);
      ASHR_i32_i32_844_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_868_inst
    process(type_cast_864_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_864_wire, type_cast_867_wire_constant, tmp_var);
      ASHR_i32_i32_868_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_894_inst
    process(type_cast_890_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_890_wire, type_cast_893_wire_constant, tmp_var);
      ASHR_i32_i32_894_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1254_inst
    process(conv153_1232, add159_1250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv153_1232, add159_1250, tmp_var);
      cmp160_1255 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1298_inst
    process(conv168_1276, add175_1294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv168_1276, add175_1294, tmp_var);
      cmp176_1299 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1804_inst
    process(conv367_1788, add373_1800) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv367_1788, add373_1800, tmp_var);
      cmp374_1805 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1847_inst
    process(conv382_1825, add389_1843) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv382_1825, add389_1843, tmp_var);
      cmp390_1848 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2368_inst
    process(conv584_2346, add591_2364) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv584_2346, add591_2364, tmp_var);
      cmp592_2369 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2412_inst
    process(conv600_2390, add607_2408) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv600_2390, add607_2408, tmp_var);
      cmp608_2413 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2930_inst
    process(conv805_2914, add811_2926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv805_2914, add811_2926, tmp_var);
      cmp812_2931 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2973_inst
    process(conv820_2951, add827_2969) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv820_2951, add827_2969, tmp_var);
      cmp828_2974 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3500_inst
    process(conv1023_3478, add1030_3496) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1023_3478, add1030_3496, tmp_var);
      cmp1031_3501 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3550_inst
    process(conv1039_3522, add1047_3546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1039_3522, add1047_3546, tmp_var);
      cmp1048_3551 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4074_inst
    process(conv1246_4058, add1252_4070) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1246_4058, add1252_4070, tmp_var);
      cmp1253_4075 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4123_inst
    process(conv1261_4095, add1269_4119) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1261_4095, add1269_4119, tmp_var);
      cmp1270_4124 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4644_inst
    process(conv1464_4622, add1471_4640) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1464_4622, add1471_4640, tmp_var);
      cmp1472_4645 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_4682_inst
    process(conv1480_4666, add1486_4678) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1480_4666, add1486_4678, tmp_var);
      cmp1487_4683 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_5200_inst
    process(conv1684_5184, add1690_5196) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1684_5184, add1690_5196, tmp_var);
      cmp1691_5201 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_5237_inst
    process(conv1699_5221, add1705_5233) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1699_5221, add1705_5233, tmp_var);
      cmp1706_5238 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1341_inst
    process(conv190_1336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv190_1336, type_cast_1340_wire_constant, tmp_var);
      div191_1342 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1890_inst
    process(conv408_1885) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv408_1885, type_cast_1889_wire_constant, tmp_var);
      div409_1891 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2455_inst
    process(conv624_2450) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv624_2450, type_cast_2454_wire_constant, tmp_var);
      div625_2456 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2468_inst
    process(conv630_2463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv630_2463, type_cast_2467_wire_constant, tmp_var);
      div631_2469 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3016_inst
    process(conv846_3011) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv846_3011, type_cast_3015_wire_constant, tmp_var);
      div847_3017 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3593_inst
    process(conv1064_3588) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1064_3588, type_cast_3592_wire_constant, tmp_var);
      div1065_3594 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3606_inst
    process(conv1070_3601) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1070_3601, type_cast_3605_wire_constant, tmp_var);
      div1071_3607 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4166_inst
    process(conv1288_4161) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1288_4161, type_cast_4165_wire_constant, tmp_var);
      div1289_4167 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4725_inst
    process(conv1503_4720) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1503_4720, type_cast_4724_wire_constant, tmp_var);
      div1504_4726 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_4744_inst
    process(mul1510_4739) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1510_4739, type_cast_4743_wire_constant, tmp_var);
      div1511_4745 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1002_inst
    process(conv69_997) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv69_997, type_cast_1001_wire_constant, tmp_var);
      div70_1003 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1244_inst
    process(conv155_1239) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1239, type_cast_1243_wire_constant, tmp_var);
      div156_1245 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1288_inst
    process(conv170_1283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv170_1283, type_cast_1287_wire_constant, tmp_var);
      div171_1289 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1514_inst
    process(conv255_1509) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv255_1509, type_cast_1513_wire_constant, tmp_var);
      div256_1515 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1837_inst
    process(conv384_1832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv384_1832, type_cast_1836_wire_constant, tmp_var);
      div385_1838 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2066_inst
    process(conv471_2061) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv471_2061, type_cast_2065_wire_constant, tmp_var);
      div472_2067 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2117_inst
    process(conv489_2112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv489_2112, type_cast_2116_wire_constant, tmp_var);
      div490_2118 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2358_inst
    process(conv586_2353) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv586_2353, type_cast_2357_wire_constant, tmp_var);
      div587_2359 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2402_inst
    process(conv602_2397) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv602_2397, type_cast_2401_wire_constant, tmp_var);
      div603_2403 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2640_inst
    process(conv693_2635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv693_2635, type_cast_2639_wire_constant, tmp_var);
      div694_2641 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2963_inst
    process(conv822_2958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv822_2958, type_cast_2962_wire_constant, tmp_var);
      div823_2964 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3198_inst
    process(mul910_3193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul910_3193, type_cast_3197_wire_constant, tmp_var);
      div911_3199 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3249_inst
    process(conv928_3244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv928_3244, type_cast_3248_wire_constant, tmp_var);
      div929_3250 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3490_inst
    process(conv1025_3485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1025_3485, type_cast_3489_wire_constant, tmp_var);
      div1026_3491 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3540_inst
    process(mul1042_3535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1042_3535, type_cast_3539_wire_constant, tmp_var);
      div1043_3541 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3784_inst
    process(mul1134_3779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1134_3779, type_cast_3783_wire_constant, tmp_var);
      div1135_3785 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4113_inst
    process(mul1264_4108) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1264_4108, type_cast_4112_wire_constant, tmp_var);
      div1265_4114 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4393_inst
    process(conv1369_4388) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1369_4388, type_cast_4392_wire_constant, tmp_var);
      div1370_4394 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_4634_inst
    process(conv1466_4629) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv1466_4629, type_cast_4633_wire_constant, tmp_var);
      div1467_4635 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_951_inst
    process(conv53_946) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv53_946, type_cast_950_wire_constant, tmp_var);
      div_952 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_4172_inst
    process(div1289_4167) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(div1289_4167, type_cast_4171_wire_constant, tmp_var);
      mul1290_4173 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_4738_inst
    process(conv1509_4733) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1509_4733, type_cast_4737_wire_constant, tmp_var);
      mul1510_4739 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1036_inst
    process(conv82_1032, conv37_831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv82_1032, conv37_831, tmp_var);
      mul83_1037 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1041_inst
    process(conv46_925, conv86_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_925, conv86_870, tmp_var);
      mul89_1042 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1095_inst
    process(sub_1091, conv31_811) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_1091, conv31_811, tmp_var);
      mul101_1096 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1105_inst
    process(sub109_1101, conv104_896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub109_1101, conv104_896, tmp_var);
      mul110_1106 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1120_inst
    process(conv60_976, conv37_831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv60_976, conv37_831, tmp_var);
      mul120_1121 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1125_inst
    process(conv46_925, conv86_870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_925, conv86_870, tmp_var);
      mul126_1126 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1414_inst
    process(conv236_1410, conv234_1395) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv236_1410, conv234_1395, tmp_var);
      mul237_1415 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1450_inst
    process(mul229_1446, conv226_1376) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul229_1446, conv226_1376, tmp_var);
      sext1719_1451 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1593_inst
    process(conv287_1589, conv234_1395) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv287_1589, conv234_1395, tmp_var);
      mul288_1594 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1598_inst
    process(conv246_1488, conv291_1434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv246_1488, conv291_1434, tmp_var);
      mul294_1599 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1651_inst
    process(sub311_1647, conv226_1376) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub311_1647, conv226_1376, tmp_var);
      mul312_1652 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1661_inst
    process(sub320_1657, conv315_1460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub320_1657, conv315_1460, tmp_var);
      mul321_1662 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1676_inst
    process(conv264_1539, conv234_1395) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv264_1539, conv234_1395, tmp_var);
      mul331_1677 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1681_inst
    process(conv246_1488, conv291_1434) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv246_1488, conv291_1434, tmp_var);
      mul337_1682 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1966_inst
    process(conv452_1962, conv450_1947) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv452_1962, conv450_1947, tmp_var);
      mul453_1967 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2002_inst
    process(mul445_1998, conv444_1932) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul445_1998, conv444_1932, tmp_var);
      sext1721_2003 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2151_inst
    process(conv504_2147, conv450_1947) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv504_2147, conv450_1947, tmp_var);
      mul505_2152 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2156_inst
    process(conv462_2040, conv508_1986) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv462_2040, conv508_1986, tmp_var);
      mul511_2157 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2209_inst
    process(sub528_2205, conv442_1928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub528_2205, conv442_1928, tmp_var);
      mul529_2210 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2219_inst
    process(sub537_2215, conv532_2012) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub537_2215, conv532_2012, tmp_var);
      mul538_2220 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2234_inst
    process(conv480_2091, conv450_1947) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv480_2091, conv450_1947, tmp_var);
      mul548_2235 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2239_inst
    process(conv462_2040, conv508_1986) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv462_2040, conv508_1986, tmp_var);
      mul554_2240 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2541_inst
    process(conv674_2537, conv672_2522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv674_2537, conv672_2522, tmp_var);
      mul675_2542 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2577_inst
    process(mul667_2573, conv666_2507) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul667_2573, conv666_2507, tmp_var);
      sext1723_2578 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2719_inst
    process(conv725_2715, conv672_2522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv725_2715, conv672_2522, tmp_var);
      mul726_2720 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2724_inst
    process(conv684_2614, conv729_2561) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv684_2614, conv729_2561, tmp_var);
      mul732_2725 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2777_inst
    process(sub749_2773, conv664_2503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub749_2773, conv664_2503, tmp_var);
      mul750_2778 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2787_inst
    process(sub758_2783, conv753_2587) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub758_2783, conv753_2587, tmp_var);
      mul759_2788 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2802_inst
    process(conv702_2665, conv672_2522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv702_2665, conv672_2522, tmp_var);
      mul769_2803 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2807_inst
    process(conv684_2614, conv729_2561) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv684_2614, conv729_2561, tmp_var);
      mul775_2808 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3092_inst
    process(conv890_3088, conv888_3073) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv890_3088, conv888_3073, tmp_var);
      mul891_3093 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3128_inst
    process(mul883_3124, conv882_3058) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul883_3124, conv882_3058, tmp_var);
      sext1725_3129 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3192_inst
    process(conv909_3187) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv909_3187, type_cast_3191_wire_constant, tmp_var);
      mul910_3193 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3283_inst
    process(conv943_3279, conv888_3073) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv943_3279, conv888_3073, tmp_var);
      mul944_3284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3288_inst
    process(conv900_3166, conv947_3112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv900_3166, conv947_3112, tmp_var);
      mul950_3289 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3341_inst
    process(sub967_3337, conv880_3054) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub967_3337, conv880_3054, tmp_var);
      mul968_3342 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3351_inst
    process(sub976_3347, conv971_3138) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub976_3347, conv971_3138, tmp_var);
      mul977_3352 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3366_inst
    process(conv919_3223, conv888_3073) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv919_3223, conv888_3073, tmp_var);
      mul987_3367 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3371_inst
    process(conv900_3166, conv947_3112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv900_3166, conv947_3112, tmp_var);
      mul993_3372 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3534_inst
    process(conv1041_3529) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1041_3529, type_cast_3533_wire_constant, tmp_var);
      mul1042_3535 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3679_inst
    process(conv1114_3675, conv1112_3660) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1114_3675, conv1112_3660, tmp_var);
      mul1115_3680 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3715_inst
    process(mul1107_3711, conv1106_3645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1107_3711, conv1106_3645, tmp_var);
      sext1727_3716 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3778_inst
    process(conv1133_3773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1133_3773, type_cast_3777_wire_constant, tmp_var);
      mul1134_3779 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3863_inst
    process(conv1166_3859, conv1112_3660) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1166_3859, conv1112_3660, tmp_var);
      mul1167_3864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3868_inst
    process(conv1124_3752, conv1170_3699) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1124_3752, conv1170_3699, tmp_var);
      mul1173_3869 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3921_inst
    process(sub1190_3917, conv1104_3641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1190_3917, conv1104_3641, tmp_var);
      mul1191_3922 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3931_inst
    process(sub1199_3927, conv1194_3725) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1199_3927, conv1194_3725, tmp_var);
      mul1200_3932 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3946_inst
    process(conv1143_3809, conv1112_3660) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1143_3809, conv1112_3660, tmp_var);
      mul1210_3947 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3951_inst
    process(conv1124_3752, conv1170_3699) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1124_3752, conv1170_3699, tmp_var);
      mul1216_3952 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4107_inst
    process(conv1263_4102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1263_4102, type_cast_4106_wire_constant, tmp_var);
      mul1264_4108 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4248_inst
    process(conv1333_4244, conv1331_4229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1333_4244, conv1331_4229, tmp_var);
      mul1334_4249 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4284_inst
    process(mul1326_4280, conv1325_4214) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1326_4280, conv1325_4214, tmp_var);
      sext1729_4285 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4427_inst
    process(conv1384_4423, conv1331_4229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1384_4423, conv1331_4229, tmp_var);
      mul1385_4428 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4432_inst
    process(conv1343_4322, conv1388_4268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1343_4322, conv1388_4268, tmp_var);
      mul1391_4433 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4485_inst
    process(sub1408_4481, conv1323_4210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1408_4481, conv1323_4210, tmp_var);
      mul1409_4486 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4495_inst
    process(sub1417_4491, conv1412_4294) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1417_4491, conv1412_4294, tmp_var);
      mul1418_4496 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4510_inst
    process(conv1360_4367, conv1331_4229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1360_4367, conv1331_4229, tmp_var);
      mul1428_4511 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4515_inst
    process(conv1343_4322, conv1388_4268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1343_4322, conv1388_4268, tmp_var);
      mul1434_4516 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4817_inst
    process(conv1554_4813, conv1552_4798) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1554_4813, conv1552_4798, tmp_var);
      mul1555_4818 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4853_inst
    process(mul1547_4849, conv1546_4783) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1547_4849, conv1546_4783, tmp_var);
      sext1731_4854 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4989_inst
    process(conv1604_4985, conv1552_4798) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1604_4985, conv1552_4798, tmp_var);
      mul1605_4990 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_4994_inst
    process(conv1564_4890, conv1608_4837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1564_4890, conv1608_4837, tmp_var);
      mul1611_4995 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5047_inst
    process(sub1628_5043, conv1544_4779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1628_5043, conv1544_4779, tmp_var);
      mul1629_5048 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5057_inst
    process(sub1637_5053, conv1632_4863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1637_5053, conv1632_4863, tmp_var);
      mul1638_5058 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5072_inst
    process(conv1581_4935, conv1552_4798) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1581_4935, conv1552_4798, tmp_var);
      mul1648_5073 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_5077_inst
    process(conv1564_4890, conv1608_4837) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1564_4890, conv1608_4837, tmp_var);
      mul1654_5078 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_850_inst
    process(conv39_846, conv37_831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv39_846, conv37_831, tmp_var);
      mul40_851 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_886_inst
    process(mul_882, conv33_815) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_882, conv33_815, tmp_var);
      sext1717_887 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1385_inst
    process(tmp213_1360) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp213_1360, type_cast_1384_wire_constant, tmp_var);
      sext1766_1386 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1400_inst
    process(tmp217_1372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp217_1372, type_cast_1399_wire_constant, tmp_var);
      sext1718_1401 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1424_inst
    process(mul237_1415) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul237_1415, type_cast_1423_wire_constant, tmp_var);
      sext1767_1425 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1439_inst
    process(conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv248_1419, type_cast_1438_wire_constant, tmp_var);
      shl372_1440 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1445_inst
    process(conv228_1380) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv228_1380, type_cast_1444_wire_constant, tmp_var);
      mul229_1446 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1937_inst
    process(tmp429_1912) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp429_1912, type_cast_1936_wire_constant, tmp_var);
      sext1768_1938 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1952_inst
    process(tmp433_1924) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp433_1924, type_cast_1951_wire_constant, tmp_var);
      sext1720_1953 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1976_inst
    process(mul453_1967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul453_1967, type_cast_1975_wire_constant, tmp_var);
      sext1769_1977 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1991_inst
    process(conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv464_1971, type_cast_1990_wire_constant, tmp_var);
      shl590_1992 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1997_inst
    process(conv442_1928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv442_1928, type_cast_1996_wire_constant, tmp_var);
      mul445_1998 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2512_inst
    process(tmp651_2487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp651_2487, type_cast_2511_wire_constant, tmp_var);
      sext1770_2513 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2527_inst
    process(tmp655_2499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp655_2499, type_cast_2526_wire_constant, tmp_var);
      sext1722_2528 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2551_inst
    process(mul675_2542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul675_2542, type_cast_2550_wire_constant, tmp_var);
      sext1771_2552 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2566_inst
    process(conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv686_2546, type_cast_2565_wire_constant, tmp_var);
      shl810_2567 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2572_inst
    process(conv664_2503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv664_2503, type_cast_2571_wire_constant, tmp_var);
      mul667_2573 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3063_inst
    process(tmp867_3038) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp867_3038, type_cast_3062_wire_constant, tmp_var);
      sext1772_3064 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3078_inst
    process(tmp871_3050) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp871_3050, type_cast_3077_wire_constant, tmp_var);
      sext1724_3079 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3102_inst
    process(mul891_3093) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul891_3093, type_cast_3101_wire_constant, tmp_var);
      sext1773_3103 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3117_inst
    process(conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv902_3097, type_cast_3116_wire_constant, tmp_var);
      shl1029_3118 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3123_inst
    process(conv880_3054) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv880_3054, type_cast_3122_wire_constant, tmp_var);
      mul883_3124 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3650_inst
    process(tmp1091_3625) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1091_3625, type_cast_3649_wire_constant, tmp_var);
      sext1774_3651 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3665_inst
    process(tmp1095_3637) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1095_3637, type_cast_3664_wire_constant, tmp_var);
      sext1726_3666 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3689_inst
    process(mul1115_3680) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1115_3680, type_cast_3688_wire_constant, tmp_var);
      sext1775_3690 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3704_inst
    process(conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1126_3684, type_cast_3703_wire_constant, tmp_var);
      shl1251_3705 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3710_inst
    process(conv1104_3641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1104_3641, type_cast_3709_wire_constant, tmp_var);
      mul1107_3711 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4219_inst
    process(tmp1310_4194) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1310_4194, type_cast_4218_wire_constant, tmp_var);
      sext1776_4220 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4234_inst
    process(tmp1314_4206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1314_4206, type_cast_4233_wire_constant, tmp_var);
      sext1728_4235 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4258_inst
    process(mul1334_4249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1334_4249, type_cast_4257_wire_constant, tmp_var);
      sext1777_4259 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4273_inst
    process(conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1345_4253, type_cast_4272_wire_constant, tmp_var);
      shl1470_4274 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4279_inst
    process(conv1323_4210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1323_4210, type_cast_4278_wire_constant, tmp_var);
      mul1326_4280 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4788_inst
    process(tmp1531_4763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1531_4763, type_cast_4787_wire_constant, tmp_var);
      sext1778_4789 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4803_inst
    process(tmp1535_4775) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp1535_4775, type_cast_4802_wire_constant, tmp_var);
      sext1730_4804 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4827_inst
    process(mul1555_4818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul1555_4818, type_cast_4826_wire_constant, tmp_var);
      sext1779_4828 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4842_inst
    process(conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1566_4822, type_cast_4841_wire_constant, tmp_var);
      shl1689_4843 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_4848_inst
    process(conv1544_4779) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1544_4779, type_cast_4847_wire_constant, tmp_var);
      mul1547_4849 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_820_inst
    process(tmp21_795) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp21_795, type_cast_819_wire_constant, tmp_var);
      sext1764_821 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_836_inst
    process(tmp24_807) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(tmp24_807, type_cast_835_wire_constant, tmp_var);
      sext_837 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_860_inst
    process(mul40_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul40_851, type_cast_859_wire_constant, tmp_var);
      sext1765_861 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_875_inst
    process(conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_855, type_cast_874_wire_constant, tmp_var);
      shl_876 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_881_inst
    process(conv31_811) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv31_811, type_cast_880_wire_constant, tmp_var);
      mul_882 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1014_inst
    process(type_cast_1011_wire, type_cast_1013_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1011_wire, type_cast_1013_wire, tmp_var);
      cmp74_1015 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1205_inst
    process(type_cast_1202_wire, type_cast_1204_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1202_wire, type_cast_1204_wire, tmp_var);
      cmp143_1206 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1494_inst
    process(type_cast_1491_wire, type_cast_1493_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1491_wire, type_cast_1493_wire, tmp_var);
      cmp249_1495 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1526_inst
    process(type_cast_1523_wire, type_cast_1525_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1523_wire, type_cast_1525_wire, tmp_var);
      cmp260_1527 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1545_inst
    process(type_cast_1542_wire, type_cast_1544_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1542_wire, type_cast_1544_wire, tmp_var);
      cmp267_1546 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1571_inst
    process(type_cast_1568_wire, type_cast_1570_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1568_wire, type_cast_1570_wire, tmp_var);
      cmp277_1572 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1761_inst
    process(type_cast_1758_wire, type_cast_1760_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1758_wire, type_cast_1760_wire, tmp_var);
      cmp356_1762 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2046_inst
    process(type_cast_2043_wire, type_cast_2045_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2043_wire, type_cast_2045_wire, tmp_var);
      cmp465_2047 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2078_inst
    process(type_cast_2075_wire, type_cast_2077_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2075_wire, type_cast_2077_wire, tmp_var);
      cmp476_2079 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2097_inst
    process(type_cast_2094_wire, type_cast_2096_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2094_wire, type_cast_2096_wire, tmp_var);
      cmp483_2098 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2129_inst
    process(type_cast_2126_wire, type_cast_2128_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2126_wire, type_cast_2128_wire, tmp_var);
      cmp494_2130 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2319_inst
    process(type_cast_2316_wire, type_cast_2318_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2316_wire, type_cast_2318_wire, tmp_var);
      cmp573_2320 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2620_inst
    process(type_cast_2617_wire, type_cast_2619_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2617_wire, type_cast_2619_wire, tmp_var);
      cmp687_2621 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2652_inst
    process(type_cast_2649_wire, type_cast_2651_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2649_wire, type_cast_2651_wire, tmp_var);
      cmp698_2653 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2671_inst
    process(type_cast_2668_wire, type_cast_2670_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2668_wire, type_cast_2670_wire, tmp_var);
      cmp705_2672 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2697_inst
    process(type_cast_2694_wire, type_cast_2696_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2694_wire, type_cast_2696_wire, tmp_var);
      cmp715_2698 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2887_inst
    process(type_cast_2884_wire, type_cast_2886_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2884_wire, type_cast_2886_wire, tmp_var);
      cmp794_2888 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3172_inst
    process(type_cast_3169_wire, type_cast_3171_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3169_wire, type_cast_3171_wire, tmp_var);
      cmp903_3173 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3210_inst
    process(type_cast_3207_wire, type_cast_3209_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3207_wire, type_cast_3209_wire, tmp_var);
      cmp915_3211 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3229_inst
    process(type_cast_3226_wire, type_cast_3228_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3226_wire, type_cast_3228_wire, tmp_var);
      cmp922_3230 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3261_inst
    process(type_cast_3258_wire, type_cast_3260_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3258_wire, type_cast_3260_wire, tmp_var);
      cmp933_3262 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3451_inst
    process(type_cast_3448_wire, type_cast_3450_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3448_wire, type_cast_3450_wire, tmp_var);
      cmp1012_3452 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3758_inst
    process(type_cast_3755_wire, type_cast_3757_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3755_wire, type_cast_3757_wire, tmp_var);
      cmp1127_3759 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3796_inst
    process(type_cast_3793_wire, type_cast_3795_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3793_wire, type_cast_3795_wire, tmp_var);
      cmp1139_3797 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3815_inst
    process(type_cast_3812_wire, type_cast_3814_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3812_wire, type_cast_3814_wire, tmp_var);
      cmp1146_3816 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3841_inst
    process(type_cast_3838_wire, type_cast_3840_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3838_wire, type_cast_3840_wire, tmp_var);
      cmp1156_3842 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4031_inst
    process(type_cast_4028_wire, type_cast_4030_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4028_wire, type_cast_4030_wire, tmp_var);
      cmp1235_4032 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4328_inst
    process(type_cast_4325_wire, type_cast_4327_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4325_wire, type_cast_4327_wire, tmp_var);
      cmp1346_4329 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4354_inst
    process(type_cast_4351_wire, type_cast_4353_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4351_wire, type_cast_4353_wire, tmp_var);
      cmp1356_4355 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4373_inst
    process(type_cast_4370_wire, type_cast_4372_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4370_wire, type_cast_4372_wire, tmp_var);
      cmp1363_4374 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4405_inst
    process(type_cast_4402_wire, type_cast_4404_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4402_wire, type_cast_4404_wire, tmp_var);
      cmp1374_4406 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4595_inst
    process(type_cast_4592_wire, type_cast_4594_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4592_wire, type_cast_4594_wire, tmp_var);
      cmp1453_4596 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4896_inst
    process(type_cast_4893_wire, type_cast_4895_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4893_wire, type_cast_4895_wire, tmp_var);
      cmp1567_4897 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4922_inst
    process(type_cast_4919_wire, type_cast_4921_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4919_wire, type_cast_4921_wire, tmp_var);
      cmp1577_4923 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4941_inst
    process(type_cast_4938_wire, type_cast_4940_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4938_wire, type_cast_4940_wire, tmp_var);
      cmp1584_4942 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_4967_inst
    process(type_cast_4964_wire, type_cast_4966_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_4964_wire, type_cast_4966_wire, tmp_var);
      cmp1594_4968 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_5157_inst
    process(type_cast_5154_wire, type_cast_5156_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_5154_wire, type_cast_5156_wire, tmp_var);
      cmp1673_5158 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_931_inst
    process(type_cast_928_wire, type_cast_930_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_928_wire, type_cast_930_wire, tmp_var);
      cmp_932 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_963_inst
    process(type_cast_960_wire, type_cast_962_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_960_wire, type_cast_962_wire, tmp_var);
      cmp56_964 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_982_inst
    process(type_cast_979_wire, type_cast_981_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_979_wire, type_cast_981_wire, tmp_var);
      cmp63_983 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1090_inst
    process(conv60_976, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv60_976, conv48_855, tmp_var);
      sub_1091 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1100_inst
    process(conv46_925, conv48_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv46_925, conv48_855, tmp_var);
      sub109_1101 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1646_inst
    process(conv264_1539, conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv264_1539, conv248_1419, tmp_var);
      sub311_1647 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1656_inst
    process(conv246_1488, conv248_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv246_1488, conv248_1419, tmp_var);
      sub320_1657 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2204_inst
    process(conv480_2091, conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv480_2091, conv464_1971, tmp_var);
      sub528_2205 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2214_inst
    process(conv462_2040, conv464_1971) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv462_2040, conv464_1971, tmp_var);
      sub537_2215 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2772_inst
    process(conv702_2665, conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv702_2665, conv686_2546, tmp_var);
      sub749_2773 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2782_inst
    process(conv684_2614, conv686_2546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv684_2614, conv686_2546, tmp_var);
      sub758_2783 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3336_inst
    process(conv919_3223, conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv919_3223, conv902_3097, tmp_var);
      sub967_3337 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3346_inst
    process(conv900_3166, conv902_3097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv900_3166, conv902_3097, tmp_var);
      sub976_3347 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3916_inst
    process(conv1143_3809, conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1143_3809, conv1126_3684, tmp_var);
      sub1190_3917 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3926_inst
    process(conv1124_3752, conv1126_3684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1124_3752, conv1126_3684, tmp_var);
      sub1199_3927 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4480_inst
    process(conv1360_4367, conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1360_4367, conv1345_4253, tmp_var);
      sub1408_4481 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_4490_inst
    process(conv1343_4322, conv1345_4253) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1343_4322, conv1345_4253, tmp_var);
      sub1417_4491 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_5042_inst
    process(conv1581_4935, conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1581_4935, conv1566_4822, tmp_var);
      sub1628_5043 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_5052_inst
    process(conv1564_4890, conv1566_4822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1564_4890, conv1566_4822, tmp_var);
      sub1637_5053 <= tmp_var; --
    end process;
    -- shared split operator group (380) : array_obj_ref_1072_index_offset 
    ApIntAdd_group_380: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1071_scaled;
      array_obj_ref_1072_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1072_index_offset_req_0;
      array_obj_ref_1072_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1072_index_offset_req_1;
      array_obj_ref_1072_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_380_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_380_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_380",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 380
    -- shared split operator group (381) : array_obj_ref_1155_index_offset 
    ApIntAdd_group_381: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom130_1154_scaled;
      array_obj_ref_1155_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1155_index_offset_req_0;
      array_obj_ref_1155_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1155_index_offset_req_1;
      array_obj_ref_1155_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_381_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_381_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_381",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 381
    -- shared split operator group (382) : array_obj_ref_1180_index_offset 
    ApIntAdd_group_382: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom135_1179_scaled;
      array_obj_ref_1180_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1180_index_offset_req_0;
      array_obj_ref_1180_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1180_index_offset_req_1;
      array_obj_ref_1180_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_382_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_382_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_382",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 382
    -- shared split operator group (383) : array_obj_ref_1628_index_offset 
    ApIntAdd_group_383: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom298_1627_scaled;
      array_obj_ref_1628_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1628_index_offset_req_0;
      array_obj_ref_1628_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1628_index_offset_req_1;
      array_obj_ref_1628_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_383_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_383_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_383",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 383
    -- shared split operator group (384) : array_obj_ref_1711_index_offset 
    ApIntAdd_group_384: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom341_1710_scaled;
      array_obj_ref_1711_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1711_index_offset_req_0;
      array_obj_ref_1711_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1711_index_offset_req_1;
      array_obj_ref_1711_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_384_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_384_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_384",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 384
    -- shared split operator group (385) : array_obj_ref_1736_index_offset 
    ApIntAdd_group_385: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom346_1735_scaled;
      array_obj_ref_1736_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1736_index_offset_req_0;
      array_obj_ref_1736_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1736_index_offset_req_1;
      array_obj_ref_1736_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_385_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_385_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_385",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 385
    -- shared split operator group (386) : array_obj_ref_2186_index_offset 
    ApIntAdd_group_386: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom515_2185_scaled;
      array_obj_ref_2186_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2186_index_offset_req_0;
      array_obj_ref_2186_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2186_index_offset_req_1;
      array_obj_ref_2186_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_386_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_386_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_386",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 386
    -- shared split operator group (387) : array_obj_ref_2269_index_offset 
    ApIntAdd_group_387: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom558_2268_scaled;
      array_obj_ref_2269_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2269_index_offset_req_0;
      array_obj_ref_2269_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2269_index_offset_req_1;
      array_obj_ref_2269_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_387_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_387_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_387",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 387
    -- shared split operator group (388) : array_obj_ref_2294_index_offset 
    ApIntAdd_group_388: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom563_2293_scaled;
      array_obj_ref_2294_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2294_index_offset_req_0;
      array_obj_ref_2294_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2294_index_offset_req_1;
      array_obj_ref_2294_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_388_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_388_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_388",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 388
    -- shared split operator group (389) : array_obj_ref_2754_index_offset 
    ApIntAdd_group_389: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom736_2753_scaled;
      array_obj_ref_2754_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2754_index_offset_req_0;
      array_obj_ref_2754_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2754_index_offset_req_1;
      array_obj_ref_2754_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_389_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_389_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_389",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 389
    -- shared split operator group (390) : array_obj_ref_2837_index_offset 
    ApIntAdd_group_390: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom779_2836_scaled;
      array_obj_ref_2837_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2837_index_offset_req_0;
      array_obj_ref_2837_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2837_index_offset_req_1;
      array_obj_ref_2837_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_390_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_390_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_390",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 390
    -- shared split operator group (391) : array_obj_ref_2862_index_offset 
    ApIntAdd_group_391: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom784_2861_scaled;
      array_obj_ref_2862_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2862_index_offset_req_0;
      array_obj_ref_2862_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2862_index_offset_req_1;
      array_obj_ref_2862_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_391_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_391_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_391",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 391
    -- shared split operator group (392) : array_obj_ref_3318_index_offset 
    ApIntAdd_group_392: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom954_3317_scaled;
      array_obj_ref_3318_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3318_index_offset_req_0;
      array_obj_ref_3318_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3318_index_offset_req_1;
      array_obj_ref_3318_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_392_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_392_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_392",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 392
    -- shared split operator group (393) : array_obj_ref_3401_index_offset 
    ApIntAdd_group_393: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom997_3400_scaled;
      array_obj_ref_3401_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3401_index_offset_req_0;
      array_obj_ref_3401_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3401_index_offset_req_1;
      array_obj_ref_3401_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_393_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_393_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_393",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 393
    -- shared split operator group (394) : array_obj_ref_3426_index_offset 
    ApIntAdd_group_394: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1002_3425_scaled;
      array_obj_ref_3426_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3426_index_offset_req_0;
      array_obj_ref_3426_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3426_index_offset_req_1;
      array_obj_ref_3426_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_394_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_394_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_394",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 394
    -- shared split operator group (395) : array_obj_ref_3898_index_offset 
    ApIntAdd_group_395: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1177_3897_scaled;
      array_obj_ref_3898_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3898_index_offset_req_0;
      array_obj_ref_3898_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3898_index_offset_req_1;
      array_obj_ref_3898_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_395_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_395_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_395",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 395
    -- shared split operator group (396) : array_obj_ref_3981_index_offset 
    ApIntAdd_group_396: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1220_3980_scaled;
      array_obj_ref_3981_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3981_index_offset_req_0;
      array_obj_ref_3981_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3981_index_offset_req_1;
      array_obj_ref_3981_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_396_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_396_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_396",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 396
    -- shared split operator group (397) : array_obj_ref_4006_index_offset 
    ApIntAdd_group_397: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1225_4005_scaled;
      array_obj_ref_4006_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4006_index_offset_req_0;
      array_obj_ref_4006_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4006_index_offset_req_1;
      array_obj_ref_4006_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_397_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_397_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_397",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 397
    -- shared split operator group (398) : array_obj_ref_4462_index_offset 
    ApIntAdd_group_398: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1395_4461_scaled;
      array_obj_ref_4462_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4462_index_offset_req_0;
      array_obj_ref_4462_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4462_index_offset_req_1;
      array_obj_ref_4462_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_398_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_398_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_398",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 398
    -- shared split operator group (399) : array_obj_ref_4545_index_offset 
    ApIntAdd_group_399: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1438_4544_scaled;
      array_obj_ref_4545_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4545_index_offset_req_0;
      array_obj_ref_4545_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4545_index_offset_req_1;
      array_obj_ref_4545_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_399_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_399_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_399",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 399
    -- shared split operator group (400) : array_obj_ref_4570_index_offset 
    ApIntAdd_group_400: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1443_4569_scaled;
      array_obj_ref_4570_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_4570_index_offset_req_0;
      array_obj_ref_4570_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_4570_index_offset_req_1;
      array_obj_ref_4570_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_400_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_400_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_400",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 400
    -- shared split operator group (401) : array_obj_ref_5024_index_offset 
    ApIntAdd_group_401: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1615_5023_scaled;
      array_obj_ref_5024_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_5024_index_offset_req_0;
      array_obj_ref_5024_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_5024_index_offset_req_1;
      array_obj_ref_5024_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_401_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_401_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_401",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 401
    -- shared split operator group (402) : array_obj_ref_5107_index_offset 
    ApIntAdd_group_402: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1658_5106_scaled;
      array_obj_ref_5107_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_5107_index_offset_req_0;
      array_obj_ref_5107_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_5107_index_offset_req_1;
      array_obj_ref_5107_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_402_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_402_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_402",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 402
    -- shared split operator group (403) : array_obj_ref_5132_index_offset 
    ApIntAdd_group_403: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1663_5131_scaled;
      array_obj_ref_5132_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_5132_index_offset_req_0;
      array_obj_ref_5132_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_5132_index_offset_req_1;
      array_obj_ref_5132_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_403_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_403_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_403",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 403
    -- unary operator type_cast_1025_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_913, tmp_var);
      type_cast_1025_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1030_inst
    process(jx_x1_899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_899, tmp_var);
      type_cast_1030_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1065_inst
    process(shr_1061) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1061, tmp_var);
      type_cast_1065_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1084_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_913, tmp_var);
      type_cast_1084_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1148_inst
    process(shr129_1145) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr129_1145, tmp_var);
      type_cast_1148_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1173_inst
    process(shr134_1170) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr134_1170, tmp_var);
      type_cast_1173_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1191_inst
    process(kx_x1_913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_913, tmp_var);
      type_cast_1191_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1230_inst
    process(inc_1227) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1227, tmp_var);
      type_cast_1230_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1274_inst
    process(inc165x_xix_x2_1264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc165x_xix_x2_1264, tmp_var);
      type_cast_1274_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1486_inst
    process(i194x_x2_1469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i194x_x2_1469, tmp_var);
      type_cast_1486_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1537_inst
    process(j240x_x1_1463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j240x_x1_1463, tmp_var);
      type_cast_1537_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1582_inst
    process(k186x_x1_1476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k186x_x1_1476, tmp_var);
      type_cast_1582_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1587_inst
    process(j240x_x1_1463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j240x_x1_1463, tmp_var);
      type_cast_1587_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1621_inst
    process(shr297_1618) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr297_1618, tmp_var);
      type_cast_1621_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1640_inst
    process(k186x_x1_1476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k186x_x1_1476, tmp_var);
      type_cast_1640_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1704_inst
    process(shr340_1701) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr340_1701, tmp_var);
      type_cast_1704_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1729_inst
    process(shr345_1726) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr345_1726, tmp_var);
      type_cast_1729_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1747_inst
    process(k186x_x1_1476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k186x_x1_1476, tmp_var);
      type_cast_1747_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1786_inst
    process(inc365_1783) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc365_1783, tmp_var);
      type_cast_1786_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1823_inst
    process(inc379x_xi194x_x2_1814) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc379x_xi194x_x2_1814, tmp_var);
      type_cast_1823_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2038_inst
    process(i406x_x2_2022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i406x_x2_2022, tmp_var);
      type_cast_2038_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2089_inst
    process(j456x_x1_2028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j456x_x1_2028, tmp_var);
      type_cast_2089_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2140_inst
    process(k402x_x1_2015) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k402x_x1_2015, tmp_var);
      type_cast_2140_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2145_inst
    process(j456x_x1_2028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j456x_x1_2028, tmp_var);
      type_cast_2145_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2179_inst
    process(shr514_2176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr514_2176, tmp_var);
      type_cast_2179_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2198_inst
    process(k402x_x1_2015) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k402x_x1_2015, tmp_var);
      type_cast_2198_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2262_inst
    process(shr557_2259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr557_2259, tmp_var);
      type_cast_2262_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2287_inst
    process(shr562_2284) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr562_2284, tmp_var);
      type_cast_2287_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2305_inst
    process(k402x_x1_2015) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k402x_x1_2015, tmp_var);
      type_cast_2305_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2344_inst
    process(inc582_2341) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc582_2341, tmp_var);
      type_cast_2344_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2388_inst
    process(inc597x_xi406x_x2_2378) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc597x_xi406x_x2_2378, tmp_var);
      type_cast_2388_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2612_inst
    process(i628x_x2_2597) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i628x_x2_2597, tmp_var);
      type_cast_2612_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2663_inst
    process(j678x_x1_2603) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j678x_x1_2603, tmp_var);
      type_cast_2663_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2708_inst
    process(k620x_x1_2590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k620x_x1_2590, tmp_var);
      type_cast_2708_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2713_inst
    process(j678x_x1_2603) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j678x_x1_2603, tmp_var);
      type_cast_2713_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2747_inst
    process(shr735_2744) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr735_2744, tmp_var);
      type_cast_2747_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2766_inst
    process(k620x_x1_2590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k620x_x1_2590, tmp_var);
      type_cast_2766_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2830_inst
    process(shr778_2827) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr778_2827, tmp_var);
      type_cast_2830_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2855_inst
    process(shr783_2852) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr783_2852, tmp_var);
      type_cast_2855_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2873_inst
    process(k620x_x1_2590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k620x_x1_2590, tmp_var);
      type_cast_2873_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2912_inst
    process(inc803_2909) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc803_2909, tmp_var);
      type_cast_2912_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2949_inst
    process(inc817x_xi628x_x2_2940) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc817x_xi628x_x2_2940, tmp_var);
      type_cast_2949_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3164_inst
    process(i844x_x2_3148) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i844x_x2_3148, tmp_var);
      type_cast_3164_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3221_inst
    process(j894x_x1_3154) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j894x_x1_3154, tmp_var);
      type_cast_3221_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3272_inst
    process(k840x_x1_3141) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k840x_x1_3141, tmp_var);
      type_cast_3272_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3277_inst
    process(j894x_x1_3154) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j894x_x1_3154, tmp_var);
      type_cast_3277_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3311_inst
    process(shr953_3308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr953_3308, tmp_var);
      type_cast_3311_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3330_inst
    process(k840x_x1_3141) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k840x_x1_3141, tmp_var);
      type_cast_3330_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3394_inst
    process(shr996_3391) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr996_3391, tmp_var);
      type_cast_3394_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3419_inst
    process(shr1001_3416) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1001_3416, tmp_var);
      type_cast_3419_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3437_inst
    process(k840x_x1_3141) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k840x_x1_3141, tmp_var);
      type_cast_3437_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3476_inst
    process(inc1021_3473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1021_3473, tmp_var);
      type_cast_3476_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3520_inst
    process(inc1036x_xi844x_x2_3510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1036x_xi844x_x2_3510, tmp_var);
      type_cast_3520_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3750_inst
    process(i1068x_x2_3735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1068x_x2_3735, tmp_var);
      type_cast_3750_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3807_inst
    process(j1118x_x1_3741) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1118x_x1_3741, tmp_var);
      type_cast_3807_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3852_inst
    process(k1060x_x1_3728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1060x_x1_3728, tmp_var);
      type_cast_3852_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3857_inst
    process(j1118x_x1_3741) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1118x_x1_3741, tmp_var);
      type_cast_3857_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3891_inst
    process(shr1176_3888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1176_3888, tmp_var);
      type_cast_3891_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3910_inst
    process(k1060x_x1_3728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1060x_x1_3728, tmp_var);
      type_cast_3910_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3974_inst
    process(shr1219_3971) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1219_3971, tmp_var);
      type_cast_3974_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3999_inst
    process(shr1224_3996) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1224_3996, tmp_var);
      type_cast_3999_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4017_inst
    process(k1060x_x1_3728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1060x_x1_3728, tmp_var);
      type_cast_4017_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4056_inst
    process(inc1244_4053) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1244_4053, tmp_var);
      type_cast_4056_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4093_inst
    process(inc1258x_xi1068x_x2_4084) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1258x_xi1068x_x2_4084, tmp_var);
      type_cast_4093_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4320_inst
    process(i1286x_x2_4304) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1286x_x2_4304, tmp_var);
      type_cast_4320_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4365_inst
    process(j1337x_x1_4310) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1337x_x1_4310, tmp_var);
      type_cast_4365_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4416_inst
    process(k1282x_x1_4297) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1282x_x1_4297, tmp_var);
      type_cast_4416_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4421_inst
    process(j1337x_x1_4310) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1337x_x1_4310, tmp_var);
      type_cast_4421_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4455_inst
    process(shr1394_4452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1394_4452, tmp_var);
      type_cast_4455_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4474_inst
    process(k1282x_x1_4297) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1282x_x1_4297, tmp_var);
      type_cast_4474_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4538_inst
    process(shr1437_4535) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1437_4535, tmp_var);
      type_cast_4538_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4563_inst
    process(shr1442_4560) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1442_4560, tmp_var);
      type_cast_4563_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4581_inst
    process(k1282x_x1_4297) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1282x_x1_4297, tmp_var);
      type_cast_4581_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4620_inst
    process(inc1462_4617) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1462_4617, tmp_var);
      type_cast_4620_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4664_inst
    process(inc1477x_xi1286x_x2_4654) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1477x_xi1286x_x2_4654, tmp_var);
      type_cast_4664_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4888_inst
    process(i1507x_x2_4873) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1507x_x2_4873, tmp_var);
      type_cast_4888_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4933_inst
    process(j1558x_x1_4879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1558x_x1_4879, tmp_var);
      type_cast_4933_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4978_inst
    process(k1499x_x1_4866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1499x_x1_4866, tmp_var);
      type_cast_4978_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_4983_inst
    process(j1558x_x1_4879) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1558x_x1_4879, tmp_var);
      type_cast_4983_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5017_inst
    process(shr1614_5014) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1614_5014, tmp_var);
      type_cast_5017_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5036_inst
    process(k1499x_x1_4866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1499x_x1_4866, tmp_var);
      type_cast_5036_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5100_inst
    process(shr1657_5097) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1657_5097, tmp_var);
      type_cast_5100_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5125_inst
    process(shr1662_5122) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1662_5122, tmp_var);
      type_cast_5125_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5143_inst
    process(k1499x_x1_4866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1499x_x1_4866, tmp_var);
      type_cast_5143_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5182_inst
    process(inc1682_5179) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1682_5179, tmp_var);
      type_cast_5182_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_5219_inst
    process(inc1696x_xi1507x_x2_5210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1696x_xi1507x_x2_5210, tmp_var);
      type_cast_5219_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_923_inst
    process(ix_x2_906) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", ix_x2_906, tmp_var);
      type_cast_923_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_974_inst
    process(jx_x1_899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_899, tmp_var);
      type_cast_974_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_col_high_4060_load_0 LOAD_col_high_1899_load_0 LOAD_col_high_1790_load_0 LOAD_col_high_782_load_0 LOAD_col_high_992_load_0 LOAD_col_high_3025_load_0 LOAD_col_high_2681_load_0 LOAD_col_high_1234_load_0 LOAD_col_high_2916_load_0 LOAD_col_high_1331_load_0 LOAD_col_high_1555_load_0 LOAD_col_high_2107_load_0 LOAD_col_high_3825_load_0 LOAD_col_high_2348_load_0 LOAD_col_high_2445_load_0 LOAD_col_high_4181_load_0 LOAD_col_high_3239_load_0 LOAD_col_high_4951_load_0 LOAD_col_high_4624_load_0 LOAD_col_high_3480_load_0 LOAD_col_high_3583_load_0 LOAD_col_high_4715_load_0 LOAD_col_high_4383_load_0 LOAD_col_high_5186_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 23 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 23 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 23 downto 0);
      signal guard_vector : std_logic_vector( 23 downto 0);
      constant inBUFs : IntegerArray(23 downto 0) := (23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(23 downto 0) := (23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(23 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false);
      constant guardBuffering: IntegerArray(23 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2);
      -- 
    begin -- 
      reqL_unguarded(23) <= LOAD_col_high_4060_load_0_req_0;
      reqL_unguarded(22) <= LOAD_col_high_1899_load_0_req_0;
      reqL_unguarded(21) <= LOAD_col_high_1790_load_0_req_0;
      reqL_unguarded(20) <= LOAD_col_high_782_load_0_req_0;
      reqL_unguarded(19) <= LOAD_col_high_992_load_0_req_0;
      reqL_unguarded(18) <= LOAD_col_high_3025_load_0_req_0;
      reqL_unguarded(17) <= LOAD_col_high_2681_load_0_req_0;
      reqL_unguarded(16) <= LOAD_col_high_1234_load_0_req_0;
      reqL_unguarded(15) <= LOAD_col_high_2916_load_0_req_0;
      reqL_unguarded(14) <= LOAD_col_high_1331_load_0_req_0;
      reqL_unguarded(13) <= LOAD_col_high_1555_load_0_req_0;
      reqL_unguarded(12) <= LOAD_col_high_2107_load_0_req_0;
      reqL_unguarded(11) <= LOAD_col_high_3825_load_0_req_0;
      reqL_unguarded(10) <= LOAD_col_high_2348_load_0_req_0;
      reqL_unguarded(9) <= LOAD_col_high_2445_load_0_req_0;
      reqL_unguarded(8) <= LOAD_col_high_4181_load_0_req_0;
      reqL_unguarded(7) <= LOAD_col_high_3239_load_0_req_0;
      reqL_unguarded(6) <= LOAD_col_high_4951_load_0_req_0;
      reqL_unguarded(5) <= LOAD_col_high_4624_load_0_req_0;
      reqL_unguarded(4) <= LOAD_col_high_3480_load_0_req_0;
      reqL_unguarded(3) <= LOAD_col_high_3583_load_0_req_0;
      reqL_unguarded(2) <= LOAD_col_high_4715_load_0_req_0;
      reqL_unguarded(1) <= LOAD_col_high_4383_load_0_req_0;
      reqL_unguarded(0) <= LOAD_col_high_5186_load_0_req_0;
      LOAD_col_high_4060_load_0_ack_0 <= ackL_unguarded(23);
      LOAD_col_high_1899_load_0_ack_0 <= ackL_unguarded(22);
      LOAD_col_high_1790_load_0_ack_0 <= ackL_unguarded(21);
      LOAD_col_high_782_load_0_ack_0 <= ackL_unguarded(20);
      LOAD_col_high_992_load_0_ack_0 <= ackL_unguarded(19);
      LOAD_col_high_3025_load_0_ack_0 <= ackL_unguarded(18);
      LOAD_col_high_2681_load_0_ack_0 <= ackL_unguarded(17);
      LOAD_col_high_1234_load_0_ack_0 <= ackL_unguarded(16);
      LOAD_col_high_2916_load_0_ack_0 <= ackL_unguarded(15);
      LOAD_col_high_1331_load_0_ack_0 <= ackL_unguarded(14);
      LOAD_col_high_1555_load_0_ack_0 <= ackL_unguarded(13);
      LOAD_col_high_2107_load_0_ack_0 <= ackL_unguarded(12);
      LOAD_col_high_3825_load_0_ack_0 <= ackL_unguarded(11);
      LOAD_col_high_2348_load_0_ack_0 <= ackL_unguarded(10);
      LOAD_col_high_2445_load_0_ack_0 <= ackL_unguarded(9);
      LOAD_col_high_4181_load_0_ack_0 <= ackL_unguarded(8);
      LOAD_col_high_3239_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_col_high_4951_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_col_high_4624_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_col_high_3480_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_col_high_3583_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_col_high_4715_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_col_high_4383_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_col_high_5186_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(23) <= LOAD_col_high_4060_load_0_req_1;
      reqR_unguarded(22) <= LOAD_col_high_1899_load_0_req_1;
      reqR_unguarded(21) <= LOAD_col_high_1790_load_0_req_1;
      reqR_unguarded(20) <= LOAD_col_high_782_load_0_req_1;
      reqR_unguarded(19) <= LOAD_col_high_992_load_0_req_1;
      reqR_unguarded(18) <= LOAD_col_high_3025_load_0_req_1;
      reqR_unguarded(17) <= LOAD_col_high_2681_load_0_req_1;
      reqR_unguarded(16) <= LOAD_col_high_1234_load_0_req_1;
      reqR_unguarded(15) <= LOAD_col_high_2916_load_0_req_1;
      reqR_unguarded(14) <= LOAD_col_high_1331_load_0_req_1;
      reqR_unguarded(13) <= LOAD_col_high_1555_load_0_req_1;
      reqR_unguarded(12) <= LOAD_col_high_2107_load_0_req_1;
      reqR_unguarded(11) <= LOAD_col_high_3825_load_0_req_1;
      reqR_unguarded(10) <= LOAD_col_high_2348_load_0_req_1;
      reqR_unguarded(9) <= LOAD_col_high_2445_load_0_req_1;
      reqR_unguarded(8) <= LOAD_col_high_4181_load_0_req_1;
      reqR_unguarded(7) <= LOAD_col_high_3239_load_0_req_1;
      reqR_unguarded(6) <= LOAD_col_high_4951_load_0_req_1;
      reqR_unguarded(5) <= LOAD_col_high_4624_load_0_req_1;
      reqR_unguarded(4) <= LOAD_col_high_3480_load_0_req_1;
      reqR_unguarded(3) <= LOAD_col_high_3583_load_0_req_1;
      reqR_unguarded(2) <= LOAD_col_high_4715_load_0_req_1;
      reqR_unguarded(1) <= LOAD_col_high_4383_load_0_req_1;
      reqR_unguarded(0) <= LOAD_col_high_5186_load_0_req_1;
      LOAD_col_high_4060_load_0_ack_1 <= ackR_unguarded(23);
      LOAD_col_high_1899_load_0_ack_1 <= ackR_unguarded(22);
      LOAD_col_high_1790_load_0_ack_1 <= ackR_unguarded(21);
      LOAD_col_high_782_load_0_ack_1 <= ackR_unguarded(20);
      LOAD_col_high_992_load_0_ack_1 <= ackR_unguarded(19);
      LOAD_col_high_3025_load_0_ack_1 <= ackR_unguarded(18);
      LOAD_col_high_2681_load_0_ack_1 <= ackR_unguarded(17);
      LOAD_col_high_1234_load_0_ack_1 <= ackR_unguarded(16);
      LOAD_col_high_2916_load_0_ack_1 <= ackR_unguarded(15);
      LOAD_col_high_1331_load_0_ack_1 <= ackR_unguarded(14);
      LOAD_col_high_1555_load_0_ack_1 <= ackR_unguarded(13);
      LOAD_col_high_2107_load_0_ack_1 <= ackR_unguarded(12);
      LOAD_col_high_3825_load_0_ack_1 <= ackR_unguarded(11);
      LOAD_col_high_2348_load_0_ack_1 <= ackR_unguarded(10);
      LOAD_col_high_2445_load_0_ack_1 <= ackR_unguarded(9);
      LOAD_col_high_4181_load_0_ack_1 <= ackR_unguarded(8);
      LOAD_col_high_3239_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_col_high_4951_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_col_high_4624_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_col_high_3480_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_col_high_3583_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_col_high_4715_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_col_high_4383_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_col_high_5186_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_16: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_17: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_17", num_slots => 1) -- 
        port map (req => reqL_unregulated(17), -- 
          ack => ackL_unregulated(17),
          regulated_req => reqL(17),
          regulated_ack => ackL(17),
          release_req => reqR(17),
          release_ack => ackR(17),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_18: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_18", num_slots => 1) -- 
        port map (req => reqL_unregulated(18), -- 
          ack => ackL_unregulated(18),
          regulated_req => reqL(18),
          regulated_ack => ackL(18),
          release_req => reqR(18),
          release_ack => ackR(18),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_19: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_19", num_slots => 1) -- 
        port map (req => reqL_unregulated(19), -- 
          ack => ackL_unregulated(19),
          regulated_req => reqL(19),
          regulated_ack => ackL(19),
          release_req => reqR(19),
          release_ack => ackR(19),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_20: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_20", num_slots => 1) -- 
        port map (req => reqL_unregulated(20), -- 
          ack => ackL_unregulated(20),
          regulated_req => reqL(20),
          regulated_ack => ackL(20),
          release_req => reqR(20),
          release_ack => ackR(20),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_21: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_21", num_slots => 1) -- 
        port map (req => reqL_unregulated(21), -- 
          ack => ackL_unregulated(21),
          regulated_req => reqL(21),
          regulated_ack => ackL(21),
          release_req => reqR(21),
          release_ack => ackR(21),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_22: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_22", num_slots => 1) -- 
        port map (req => reqL_unregulated(22), -- 
          ack => ackL_unregulated(22),
          regulated_req => reqL(22),
          regulated_ack => ackL(22),
          release_req => reqR(22),
          release_ack => ackR(22),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_23: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_23", num_slots => 1) -- 
        port map (req => reqL_unregulated(23), -- 
          ack => ackL_unregulated(23),
          regulated_req => reqL(23),
          regulated_ack => ackL(23),
          release_req => reqR(23),
          release_ack => ackR(23),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 24, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_col_high_4060_word_address_0 & LOAD_col_high_1899_word_address_0 & LOAD_col_high_1790_word_address_0 & LOAD_col_high_782_word_address_0 & LOAD_col_high_992_word_address_0 & LOAD_col_high_3025_word_address_0 & LOAD_col_high_2681_word_address_0 & LOAD_col_high_1234_word_address_0 & LOAD_col_high_2916_word_address_0 & LOAD_col_high_1331_word_address_0 & LOAD_col_high_1555_word_address_0 & LOAD_col_high_2107_word_address_0 & LOAD_col_high_3825_word_address_0 & LOAD_col_high_2348_word_address_0 & LOAD_col_high_2445_word_address_0 & LOAD_col_high_4181_word_address_0 & LOAD_col_high_3239_word_address_0 & LOAD_col_high_4951_word_address_0 & LOAD_col_high_4624_word_address_0 & LOAD_col_high_3480_word_address_0 & LOAD_col_high_3583_word_address_0 & LOAD_col_high_4715_word_address_0 & LOAD_col_high_4383_word_address_0 & LOAD_col_high_5186_word_address_0;
      LOAD_col_high_4060_data_0 <= data_out(191 downto 184);
      LOAD_col_high_1899_data_0 <= data_out(183 downto 176);
      LOAD_col_high_1790_data_0 <= data_out(175 downto 168);
      LOAD_col_high_782_data_0 <= data_out(167 downto 160);
      LOAD_col_high_992_data_0 <= data_out(159 downto 152);
      LOAD_col_high_3025_data_0 <= data_out(151 downto 144);
      LOAD_col_high_2681_data_0 <= data_out(143 downto 136);
      LOAD_col_high_1234_data_0 <= data_out(135 downto 128);
      LOAD_col_high_2916_data_0 <= data_out(127 downto 120);
      LOAD_col_high_1331_data_0 <= data_out(119 downto 112);
      LOAD_col_high_1555_data_0 <= data_out(111 downto 104);
      LOAD_col_high_2107_data_0 <= data_out(103 downto 96);
      LOAD_col_high_3825_data_0 <= data_out(95 downto 88);
      LOAD_col_high_2348_data_0 <= data_out(87 downto 80);
      LOAD_col_high_2445_data_0 <= data_out(79 downto 72);
      LOAD_col_high_4181_data_0 <= data_out(71 downto 64);
      LOAD_col_high_3239_data_0 <= data_out(63 downto 56);
      LOAD_col_high_4951_data_0 <= data_out(55 downto 48);
      LOAD_col_high_4624_data_0 <= data_out(47 downto 40);
      LOAD_col_high_3480_data_0 <= data_out(39 downto 32);
      LOAD_col_high_3583_data_0 <= data_out(31 downto 24);
      LOAD_col_high_4715_data_0 <= data_out(23 downto 16);
      LOAD_col_high_4383_data_0 <= data_out(15 downto 8);
      LOAD_col_high_5186_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 24,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 24,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : LOAD_depth_high_1896_load_0 LOAD_depth_high_3022_load_0 LOAD_depth_high_779_load_0 LOAD_depth_high_1347_load_0 LOAD_depth_high_2474_load_0 LOAD_depth_high_4750_load_0 LOAD_depth_high_4178_load_0 LOAD_depth_high_3612_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_depth_high_1896_load_0_req_0;
      reqL_unguarded(6) <= LOAD_depth_high_3022_load_0_req_0;
      reqL_unguarded(5) <= LOAD_depth_high_779_load_0_req_0;
      reqL_unguarded(4) <= LOAD_depth_high_1347_load_0_req_0;
      reqL_unguarded(3) <= LOAD_depth_high_2474_load_0_req_0;
      reqL_unguarded(2) <= LOAD_depth_high_4750_load_0_req_0;
      reqL_unguarded(1) <= LOAD_depth_high_4178_load_0_req_0;
      reqL_unguarded(0) <= LOAD_depth_high_3612_load_0_req_0;
      LOAD_depth_high_1896_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_depth_high_3022_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_depth_high_779_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_depth_high_1347_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_depth_high_2474_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_depth_high_4750_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_depth_high_4178_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_depth_high_3612_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_depth_high_1896_load_0_req_1;
      reqR_unguarded(6) <= LOAD_depth_high_3022_load_0_req_1;
      reqR_unguarded(5) <= LOAD_depth_high_779_load_0_req_1;
      reqR_unguarded(4) <= LOAD_depth_high_1347_load_0_req_1;
      reqR_unguarded(3) <= LOAD_depth_high_2474_load_0_req_1;
      reqR_unguarded(2) <= LOAD_depth_high_4750_load_0_req_1;
      reqR_unguarded(1) <= LOAD_depth_high_4178_load_0_req_1;
      reqR_unguarded(0) <= LOAD_depth_high_3612_load_0_req_1;
      LOAD_depth_high_1896_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_depth_high_3022_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_depth_high_779_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_depth_high_1347_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_depth_high_2474_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_depth_high_4750_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_depth_high_4178_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_depth_high_3612_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_depth_high_1896_word_address_0 & LOAD_depth_high_3022_word_address_0 & LOAD_depth_high_779_word_address_0 & LOAD_depth_high_1347_word_address_0 & LOAD_depth_high_2474_word_address_0 & LOAD_depth_high_4750_word_address_0 & LOAD_depth_high_4178_word_address_0 & LOAD_depth_high_3612_word_address_0;
      LOAD_depth_high_1896_data_0 <= data_out(63 downto 56);
      LOAD_depth_high_3022_data_0 <= data_out(55 downto 48);
      LOAD_depth_high_779_data_0 <= data_out(47 downto 40);
      LOAD_depth_high_1347_data_0 <= data_out(39 downto 32);
      LOAD_depth_high_2474_data_0 <= data_out(31 downto 24);
      LOAD_depth_high_4750_data_0 <= data_out(23 downto 16);
      LOAD_depth_high_4178_data_0 <= data_out(15 downto 8);
      LOAD_depth_high_3612_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(7 downto 0),
          mtag => memory_space_4_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : LOAD_pad_1893_load_0 LOAD_pad_776_load_0 LOAD_pad_3019_load_0 LOAD_pad_1344_load_0 LOAD_pad_2471_load_0 LOAD_pad_4175_load_0 LOAD_pad_4747_load_0 LOAD_pad_3609_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_pad_1893_load_0_req_0;
      reqL_unguarded(6) <= LOAD_pad_776_load_0_req_0;
      reqL_unguarded(5) <= LOAD_pad_3019_load_0_req_0;
      reqL_unguarded(4) <= LOAD_pad_1344_load_0_req_0;
      reqL_unguarded(3) <= LOAD_pad_2471_load_0_req_0;
      reqL_unguarded(2) <= LOAD_pad_4175_load_0_req_0;
      reqL_unguarded(1) <= LOAD_pad_4747_load_0_req_0;
      reqL_unguarded(0) <= LOAD_pad_3609_load_0_req_0;
      LOAD_pad_1893_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_pad_776_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_pad_3019_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_pad_1344_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_pad_2471_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_pad_4175_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_pad_4747_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_pad_3609_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_pad_1893_load_0_req_1;
      reqR_unguarded(6) <= LOAD_pad_776_load_0_req_1;
      reqR_unguarded(5) <= LOAD_pad_3019_load_0_req_1;
      reqR_unguarded(4) <= LOAD_pad_1344_load_0_req_1;
      reqR_unguarded(3) <= LOAD_pad_2471_load_0_req_1;
      reqR_unguarded(2) <= LOAD_pad_4175_load_0_req_1;
      reqR_unguarded(1) <= LOAD_pad_4747_load_0_req_1;
      reqR_unguarded(0) <= LOAD_pad_3609_load_0_req_1;
      LOAD_pad_1893_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_pad_776_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_pad_3019_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_pad_1344_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_pad_2471_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_pad_4175_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_pad_4747_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_pad_3609_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_1893_word_address_0 & LOAD_pad_776_word_address_0 & LOAD_pad_3019_word_address_0 & LOAD_pad_1344_word_address_0 & LOAD_pad_2471_word_address_0 & LOAD_pad_4175_word_address_0 & LOAD_pad_4747_word_address_0 & LOAD_pad_3609_word_address_0;
      LOAD_pad_1893_data_0 <= data_out(63 downto 56);
      LOAD_pad_776_data_0 <= data_out(55 downto 48);
      LOAD_pad_3019_data_0 <= data_out(47 downto 40);
      LOAD_pad_1344_data_0 <= data_out(39 downto 32);
      LOAD_pad_2471_data_0 <= data_out(31 downto 24);
      LOAD_pad_4175_data_0 <= data_out(23 downto 16);
      LOAD_pad_4747_data_0 <= data_out(15 downto 8);
      LOAD_pad_3609_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : LOAD_row_high_1880_load_0 LOAD_row_high_1827_load_0 LOAD_row_high_2630_load_0 LOAD_row_high_941_load_0 LOAD_row_high_2953_load_0 LOAD_row_high_4728_load_0 LOAD_row_high_3006_load_0 LOAD_row_high_4097_load_0 LOAD_row_high_1278_load_0 LOAD_row_high_1504_load_0 LOAD_row_high_2056_load_0 LOAD_row_high_3768_load_0 LOAD_row_high_2392_load_0 LOAD_row_high_2458_load_0 LOAD_row_high_3182_load_0 LOAD_row_high_4156_load_0 LOAD_row_high_4668_load_0 LOAD_row_high_3524_load_0 LOAD_row_high_3596_load_0 LOAD_row_high_4906_load_0 LOAD_row_high_4338_load_0 LOAD_row_high_5223_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(175 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 21 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 21 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 21 downto 0);
      signal guard_vector : std_logic_vector( 21 downto 0);
      constant inBUFs : IntegerArray(21 downto 0) := (21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(21 downto 0) := (21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(21 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false);
      constant guardBuffering: IntegerArray(21 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2);
      -- 
    begin -- 
      reqL_unguarded(21) <= LOAD_row_high_1880_load_0_req_0;
      reqL_unguarded(20) <= LOAD_row_high_1827_load_0_req_0;
      reqL_unguarded(19) <= LOAD_row_high_2630_load_0_req_0;
      reqL_unguarded(18) <= LOAD_row_high_941_load_0_req_0;
      reqL_unguarded(17) <= LOAD_row_high_2953_load_0_req_0;
      reqL_unguarded(16) <= LOAD_row_high_4728_load_0_req_0;
      reqL_unguarded(15) <= LOAD_row_high_3006_load_0_req_0;
      reqL_unguarded(14) <= LOAD_row_high_4097_load_0_req_0;
      reqL_unguarded(13) <= LOAD_row_high_1278_load_0_req_0;
      reqL_unguarded(12) <= LOAD_row_high_1504_load_0_req_0;
      reqL_unguarded(11) <= LOAD_row_high_2056_load_0_req_0;
      reqL_unguarded(10) <= LOAD_row_high_3768_load_0_req_0;
      reqL_unguarded(9) <= LOAD_row_high_2392_load_0_req_0;
      reqL_unguarded(8) <= LOAD_row_high_2458_load_0_req_0;
      reqL_unguarded(7) <= LOAD_row_high_3182_load_0_req_0;
      reqL_unguarded(6) <= LOAD_row_high_4156_load_0_req_0;
      reqL_unguarded(5) <= LOAD_row_high_4668_load_0_req_0;
      reqL_unguarded(4) <= LOAD_row_high_3524_load_0_req_0;
      reqL_unguarded(3) <= LOAD_row_high_3596_load_0_req_0;
      reqL_unguarded(2) <= LOAD_row_high_4906_load_0_req_0;
      reqL_unguarded(1) <= LOAD_row_high_4338_load_0_req_0;
      reqL_unguarded(0) <= LOAD_row_high_5223_load_0_req_0;
      LOAD_row_high_1880_load_0_ack_0 <= ackL_unguarded(21);
      LOAD_row_high_1827_load_0_ack_0 <= ackL_unguarded(20);
      LOAD_row_high_2630_load_0_ack_0 <= ackL_unguarded(19);
      LOAD_row_high_941_load_0_ack_0 <= ackL_unguarded(18);
      LOAD_row_high_2953_load_0_ack_0 <= ackL_unguarded(17);
      LOAD_row_high_4728_load_0_ack_0 <= ackL_unguarded(16);
      LOAD_row_high_3006_load_0_ack_0 <= ackL_unguarded(15);
      LOAD_row_high_4097_load_0_ack_0 <= ackL_unguarded(14);
      LOAD_row_high_1278_load_0_ack_0 <= ackL_unguarded(13);
      LOAD_row_high_1504_load_0_ack_0 <= ackL_unguarded(12);
      LOAD_row_high_2056_load_0_ack_0 <= ackL_unguarded(11);
      LOAD_row_high_3768_load_0_ack_0 <= ackL_unguarded(10);
      LOAD_row_high_2392_load_0_ack_0 <= ackL_unguarded(9);
      LOAD_row_high_2458_load_0_ack_0 <= ackL_unguarded(8);
      LOAD_row_high_3182_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_row_high_4156_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_row_high_4668_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_row_high_3524_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_row_high_3596_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_row_high_4906_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_row_high_4338_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_row_high_5223_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(21) <= LOAD_row_high_1880_load_0_req_1;
      reqR_unguarded(20) <= LOAD_row_high_1827_load_0_req_1;
      reqR_unguarded(19) <= LOAD_row_high_2630_load_0_req_1;
      reqR_unguarded(18) <= LOAD_row_high_941_load_0_req_1;
      reqR_unguarded(17) <= LOAD_row_high_2953_load_0_req_1;
      reqR_unguarded(16) <= LOAD_row_high_4728_load_0_req_1;
      reqR_unguarded(15) <= LOAD_row_high_3006_load_0_req_1;
      reqR_unguarded(14) <= LOAD_row_high_4097_load_0_req_1;
      reqR_unguarded(13) <= LOAD_row_high_1278_load_0_req_1;
      reqR_unguarded(12) <= LOAD_row_high_1504_load_0_req_1;
      reqR_unguarded(11) <= LOAD_row_high_2056_load_0_req_1;
      reqR_unguarded(10) <= LOAD_row_high_3768_load_0_req_1;
      reqR_unguarded(9) <= LOAD_row_high_2392_load_0_req_1;
      reqR_unguarded(8) <= LOAD_row_high_2458_load_0_req_1;
      reqR_unguarded(7) <= LOAD_row_high_3182_load_0_req_1;
      reqR_unguarded(6) <= LOAD_row_high_4156_load_0_req_1;
      reqR_unguarded(5) <= LOAD_row_high_4668_load_0_req_1;
      reqR_unguarded(4) <= LOAD_row_high_3524_load_0_req_1;
      reqR_unguarded(3) <= LOAD_row_high_3596_load_0_req_1;
      reqR_unguarded(2) <= LOAD_row_high_4906_load_0_req_1;
      reqR_unguarded(1) <= LOAD_row_high_4338_load_0_req_1;
      reqR_unguarded(0) <= LOAD_row_high_5223_load_0_req_1;
      LOAD_row_high_1880_load_0_ack_1 <= ackR_unguarded(21);
      LOAD_row_high_1827_load_0_ack_1 <= ackR_unguarded(20);
      LOAD_row_high_2630_load_0_ack_1 <= ackR_unguarded(19);
      LOAD_row_high_941_load_0_ack_1 <= ackR_unguarded(18);
      LOAD_row_high_2953_load_0_ack_1 <= ackR_unguarded(17);
      LOAD_row_high_4728_load_0_ack_1 <= ackR_unguarded(16);
      LOAD_row_high_3006_load_0_ack_1 <= ackR_unguarded(15);
      LOAD_row_high_4097_load_0_ack_1 <= ackR_unguarded(14);
      LOAD_row_high_1278_load_0_ack_1 <= ackR_unguarded(13);
      LOAD_row_high_1504_load_0_ack_1 <= ackR_unguarded(12);
      LOAD_row_high_2056_load_0_ack_1 <= ackR_unguarded(11);
      LOAD_row_high_3768_load_0_ack_1 <= ackR_unguarded(10);
      LOAD_row_high_2392_load_0_ack_1 <= ackR_unguarded(9);
      LOAD_row_high_2458_load_0_ack_1 <= ackR_unguarded(8);
      LOAD_row_high_3182_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_row_high_4156_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_row_high_4668_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_row_high_3524_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_row_high_3596_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_row_high_4906_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_row_high_4338_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_row_high_5223_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_16: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_17: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_17", num_slots => 1) -- 
        port map (req => reqL_unregulated(17), -- 
          ack => ackL_unregulated(17),
          regulated_req => reqL(17),
          regulated_ack => ackL(17),
          release_req => reqR(17),
          release_ack => ackR(17),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_18: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_18", num_slots => 1) -- 
        port map (req => reqL_unregulated(18), -- 
          ack => ackL_unregulated(18),
          regulated_req => reqL(18),
          regulated_ack => ackL(18),
          release_req => reqR(18),
          release_ack => ackR(18),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_19: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_19", num_slots => 1) -- 
        port map (req => reqL_unregulated(19), -- 
          ack => ackL_unregulated(19),
          regulated_req => reqL(19),
          regulated_ack => ackL(19),
          release_req => reqR(19),
          release_ack => ackR(19),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_20: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_20", num_slots => 1) -- 
        port map (req => reqL_unregulated(20), -- 
          ack => ackL_unregulated(20),
          regulated_req => reqL(20),
          regulated_ack => ackL(20),
          release_req => reqR(20),
          release_ack => ackR(20),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_21: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_21", num_slots => 1) -- 
        port map (req => reqL_unregulated(21), -- 
          ack => ackL_unregulated(21),
          regulated_req => reqL(21),
          regulated_ack => ackL(21),
          release_req => reqR(21),
          release_ack => ackR(21),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 22, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_row_high_1880_word_address_0 & LOAD_row_high_1827_word_address_0 & LOAD_row_high_2630_word_address_0 & LOAD_row_high_941_word_address_0 & LOAD_row_high_2953_word_address_0 & LOAD_row_high_4728_word_address_0 & LOAD_row_high_3006_word_address_0 & LOAD_row_high_4097_word_address_0 & LOAD_row_high_1278_word_address_0 & LOAD_row_high_1504_word_address_0 & LOAD_row_high_2056_word_address_0 & LOAD_row_high_3768_word_address_0 & LOAD_row_high_2392_word_address_0 & LOAD_row_high_2458_word_address_0 & LOAD_row_high_3182_word_address_0 & LOAD_row_high_4156_word_address_0 & LOAD_row_high_4668_word_address_0 & LOAD_row_high_3524_word_address_0 & LOAD_row_high_3596_word_address_0 & LOAD_row_high_4906_word_address_0 & LOAD_row_high_4338_word_address_0 & LOAD_row_high_5223_word_address_0;
      LOAD_row_high_1880_data_0 <= data_out(175 downto 168);
      LOAD_row_high_1827_data_0 <= data_out(167 downto 160);
      LOAD_row_high_2630_data_0 <= data_out(159 downto 152);
      LOAD_row_high_941_data_0 <= data_out(151 downto 144);
      LOAD_row_high_2953_data_0 <= data_out(143 downto 136);
      LOAD_row_high_4728_data_0 <= data_out(135 downto 128);
      LOAD_row_high_3006_data_0 <= data_out(127 downto 120);
      LOAD_row_high_4097_data_0 <= data_out(119 downto 112);
      LOAD_row_high_1278_data_0 <= data_out(111 downto 104);
      LOAD_row_high_1504_data_0 <= data_out(103 downto 96);
      LOAD_row_high_2056_data_0 <= data_out(95 downto 88);
      LOAD_row_high_3768_data_0 <= data_out(87 downto 80);
      LOAD_row_high_2392_data_0 <= data_out(79 downto 72);
      LOAD_row_high_2458_data_0 <= data_out(71 downto 64);
      LOAD_row_high_3182_data_0 <= data_out(63 downto 56);
      LOAD_row_high_4156_data_0 <= data_out(55 downto 48);
      LOAD_row_high_4668_data_0 <= data_out(47 downto 40);
      LOAD_row_high_3524_data_0 <= data_out(39 downto 32);
      LOAD_row_high_3596_data_0 <= data_out(31 downto 24);
      LOAD_row_high_4906_data_0 <= data_out(23 downto 16);
      LOAD_row_high_4338_data_0 <= data_out(15 downto 8);
      LOAD_row_high_5223_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 1,
        num_reqs => 22,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 8,
        num_reqs => 22,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1160_load_0 ptr_deref_2842_load_0 ptr_deref_1716_load_0 ptr_deref_2274_load_0 ptr_deref_3986_load_0 ptr_deref_3406_load_0 ptr_deref_5112_load_0 ptr_deref_4550_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_1160_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2842_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_1716_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_2274_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_3986_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3406_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_5112_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4550_load_0_req_0;
      ptr_deref_1160_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2842_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_1716_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_2274_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_3986_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3406_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_5112_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4550_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_1160_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2842_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_1716_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_2274_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_3986_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3406_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_5112_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4550_load_0_req_1;
      ptr_deref_1160_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2842_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_1716_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_2274_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_3986_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3406_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_5112_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4550_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1160_word_address_0 & ptr_deref_2842_word_address_0 & ptr_deref_1716_word_address_0 & ptr_deref_2274_word_address_0 & ptr_deref_3986_word_address_0 & ptr_deref_3406_word_address_0 & ptr_deref_5112_word_address_0 & ptr_deref_4550_word_address_0;
      ptr_deref_1160_data_0 <= data_out(511 downto 448);
      ptr_deref_2842_data_0 <= data_out(447 downto 384);
      ptr_deref_1716_data_0 <= data_out(383 downto 320);
      ptr_deref_2274_data_0 <= data_out(319 downto 256);
      ptr_deref_3986_data_0 <= data_out(255 downto 192);
      ptr_deref_3406_data_0 <= data_out(191 downto 128);
      ptr_deref_5112_data_0 <= data_out(127 downto 64);
      ptr_deref_4550_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 14,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 64,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_806_load_0 ptr_deref_794_load_0 ptr_deref_1911_load_0 ptr_deref_1923_load_0 ptr_deref_3049_load_0 ptr_deref_1359_load_0 ptr_deref_1371_load_0 ptr_deref_3037_load_0 ptr_deref_2486_load_0 ptr_deref_2498_load_0 ptr_deref_3636_load_0 ptr_deref_4193_load_0 ptr_deref_4205_load_0 ptr_deref_3624_load_0 ptr_deref_4774_load_0 ptr_deref_4762_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_806_load_0_req_0;
      reqL_unguarded(14) <= ptr_deref_794_load_0_req_0;
      reqL_unguarded(13) <= ptr_deref_1911_load_0_req_0;
      reqL_unguarded(12) <= ptr_deref_1923_load_0_req_0;
      reqL_unguarded(11) <= ptr_deref_3049_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_1359_load_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1371_load_0_req_0;
      reqL_unguarded(8) <= ptr_deref_3037_load_0_req_0;
      reqL_unguarded(7) <= ptr_deref_2486_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2498_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_3636_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_4193_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_4205_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_3624_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_4774_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4762_load_0_req_0;
      ptr_deref_806_load_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_794_load_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_1911_load_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_1923_load_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_3049_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_1359_load_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1371_load_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_3037_load_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_2486_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2498_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_3636_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_4193_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_4205_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_3624_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_4774_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4762_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_806_load_0_req_1;
      reqR_unguarded(14) <= ptr_deref_794_load_0_req_1;
      reqR_unguarded(13) <= ptr_deref_1911_load_0_req_1;
      reqR_unguarded(12) <= ptr_deref_1923_load_0_req_1;
      reqR_unguarded(11) <= ptr_deref_3049_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_1359_load_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1371_load_0_req_1;
      reqR_unguarded(8) <= ptr_deref_3037_load_0_req_1;
      reqR_unguarded(7) <= ptr_deref_2486_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2498_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_3636_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_4193_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_4205_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_3624_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_4774_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4762_load_0_req_1;
      ptr_deref_806_load_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_794_load_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_1911_load_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_1923_load_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_3049_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_1359_load_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1371_load_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_3037_load_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_2486_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2498_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_3636_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_4193_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_4205_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_3624_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_4774_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4762_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup5_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup5_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup5_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_806_word_address_0 & ptr_deref_794_word_address_0 & ptr_deref_1911_word_address_0 & ptr_deref_1923_word_address_0 & ptr_deref_3049_word_address_0 & ptr_deref_1359_word_address_0 & ptr_deref_1371_word_address_0 & ptr_deref_3037_word_address_0 & ptr_deref_2486_word_address_0 & ptr_deref_2498_word_address_0 & ptr_deref_3636_word_address_0 & ptr_deref_4193_word_address_0 & ptr_deref_4205_word_address_0 & ptr_deref_3624_word_address_0 & ptr_deref_4774_word_address_0 & ptr_deref_4762_word_address_0;
      ptr_deref_806_data_0 <= data_out(511 downto 480);
      ptr_deref_794_data_0 <= data_out(479 downto 448);
      ptr_deref_1911_data_0 <= data_out(447 downto 416);
      ptr_deref_1923_data_0 <= data_out(415 downto 384);
      ptr_deref_3049_data_0 <= data_out(383 downto 352);
      ptr_deref_1359_data_0 <= data_out(351 downto 320);
      ptr_deref_1371_data_0 <= data_out(319 downto 288);
      ptr_deref_3037_data_0 <= data_out(287 downto 256);
      ptr_deref_2486_data_0 <= data_out(255 downto 224);
      ptr_deref_2498_data_0 <= data_out(223 downto 192);
      ptr_deref_3636_data_0 <= data_out(191 downto 160);
      ptr_deref_4193_data_0 <= data_out(159 downto 128);
      ptr_deref_4205_data_0 <= data_out(127 downto 96);
      ptr_deref_3624_data_0 <= data_out(95 downto 64);
      ptr_deref_4774_data_0 <= data_out(63 downto 32);
      ptr_deref_4762_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 7,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(6 downto 0),
          mtag => memory_space_6_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 32,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_727_load_0 ptr_deref_746_load_0 ptr_deref_765_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_727_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_746_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_765_load_0_req_0;
      ptr_deref_727_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_746_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_765_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_727_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_746_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_765_load_0_req_1;
      ptr_deref_727_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_746_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_765_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup6_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup6_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup6_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup6_gI: SplitGuardInterface generic map(name => "LoadGroup6_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_727_word_address_0 & ptr_deref_746_word_address_0 & ptr_deref_765_word_address_0;
      ptr_deref_727_data_0 <= data_out(95 downto 64);
      ptr_deref_746_data_0 <= data_out(63 downto 32);
      ptr_deref_765_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup6", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(6 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup6 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared store operator group (0) : STORE_col_high_752_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_col_high_752_store_0_req_0;
      STORE_col_high_752_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_col_high_752_store_0_req_1;
      STORE_col_high_752_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_col_high_752_word_address_0;
      data_in <= STORE_col_high_752_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : STORE_depth_high_771_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_depth_high_771_store_0_req_0;
      STORE_depth_high_771_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_depth_high_771_store_0_req_1;
      STORE_depth_high_771_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_depth_high_771_word_address_0;
      data_in <= STORE_depth_high_771_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : STORE_row_high_733_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_row_high_733_store_0_req_0;
      STORE_row_high_733_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_row_high_733_store_0_req_1;
      STORE_row_high_733_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_row_high_733_word_address_0;
      data_in <= STORE_row_high_733_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_3902_store_0 ptr_deref_1076_store_0 ptr_deref_2758_store_0 ptr_deref_1184_store_0 ptr_deref_4010_store_0 ptr_deref_2866_store_0 ptr_deref_1632_store_0 ptr_deref_1740_store_0 ptr_deref_2190_store_0 ptr_deref_2298_store_0 ptr_deref_5136_store_0 ptr_deref_3322_store_0 ptr_deref_3430_store_0 ptr_deref_5028_store_0 ptr_deref_4466_store_0 ptr_deref_4574_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(223 downto 0);
      signal data_in: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_3902_store_0_req_0;
      reqL_unguarded(14) <= ptr_deref_1076_store_0_req_0;
      reqL_unguarded(13) <= ptr_deref_2758_store_0_req_0;
      reqL_unguarded(12) <= ptr_deref_1184_store_0_req_0;
      reqL_unguarded(11) <= ptr_deref_4010_store_0_req_0;
      reqL_unguarded(10) <= ptr_deref_2866_store_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1632_store_0_req_0;
      reqL_unguarded(8) <= ptr_deref_1740_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_2190_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2298_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_5136_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_3322_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_3430_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_5028_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_4466_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_4574_store_0_req_0;
      ptr_deref_3902_store_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_1076_store_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_2758_store_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_1184_store_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_4010_store_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_2866_store_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1632_store_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_1740_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_2190_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2298_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_5136_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_3322_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_3430_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_5028_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_4466_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_4574_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_3902_store_0_req_1;
      reqR_unguarded(14) <= ptr_deref_1076_store_0_req_1;
      reqR_unguarded(13) <= ptr_deref_2758_store_0_req_1;
      reqR_unguarded(12) <= ptr_deref_1184_store_0_req_1;
      reqR_unguarded(11) <= ptr_deref_4010_store_0_req_1;
      reqR_unguarded(10) <= ptr_deref_2866_store_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1632_store_0_req_1;
      reqR_unguarded(8) <= ptr_deref_1740_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_2190_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2298_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_5136_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_3322_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_3430_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_5028_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_4466_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_4574_store_0_req_1;
      ptr_deref_3902_store_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_1076_store_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_2758_store_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_1184_store_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_4010_store_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_2866_store_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1632_store_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_1740_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_2190_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2298_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_5136_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_3322_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_3430_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_5028_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_4466_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_4574_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_13: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_14: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_15: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3902_word_address_0 & ptr_deref_1076_word_address_0 & ptr_deref_2758_word_address_0 & ptr_deref_1184_word_address_0 & ptr_deref_4010_word_address_0 & ptr_deref_2866_word_address_0 & ptr_deref_1632_word_address_0 & ptr_deref_1740_word_address_0 & ptr_deref_2190_word_address_0 & ptr_deref_2298_word_address_0 & ptr_deref_5136_word_address_0 & ptr_deref_3322_word_address_0 & ptr_deref_3430_word_address_0 & ptr_deref_5028_word_address_0 & ptr_deref_4466_word_address_0 & ptr_deref_4574_word_address_0;
      data_in <= ptr_deref_3902_data_0 & ptr_deref_1076_data_0 & ptr_deref_2758_data_0 & ptr_deref_1184_data_0 & ptr_deref_4010_data_0 & ptr_deref_2866_data_0 & ptr_deref_1632_data_0 & ptr_deref_1740_data_0 & ptr_deref_2190_data_0 & ptr_deref_2298_data_0 & ptr_deref_5136_data_0 & ptr_deref_3322_data_0 & ptr_deref_3430_data_0 & ptr_deref_5028_data_0 & ptr_deref_4466_data_0 & ptr_deref_4574_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 16,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared call operator group (0) : call_stmt_5270_call 
    sendOutput_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_5270_call_req_0;
      call_stmt_5270_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_5270_call_req_1;
      call_stmt_5270_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_0_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_716_call 
    testConfigure_call_group_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_716_call_req_0;
      call_stmt_716_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_716_call_req_1;
      call_stmt_716_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_1_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_716 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(43 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(9 downto 0);
  -- interface signals to connect to memory space memory_space_3
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(1 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(41 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(7 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(1 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(43 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(9 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(4 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(21 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(4 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(13 downto 7),
      memory_space_6_lr_tag => memory_space_6_lr_tag(43 downto 22),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(9 downto 5),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(13 downto 7),
      memory_space_5_lr_tag => memory_space_5_lr_tag(37 downto 19),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 32),
      memory_space_5_lc_tag => memory_space_5_lc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(1 downto 1),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 8),
      memory_space_2_sr_tag => memory_space_2_sr_tag(43 downto 22),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(9 downto 5),
      memory_space_4_sr_req => memory_space_4_sr_req(1 downto 1),
      memory_space_4_sr_ack => memory_space_4_sr_ack(1 downto 1),
      memory_space_4_sr_addr => memory_space_4_sr_addr(1 downto 1),
      memory_space_4_sr_data => memory_space_4_sr_data(15 downto 8),
      memory_space_4_sr_tag => memory_space_4_sr_tag(41 downto 21),
      memory_space_4_sc_req => memory_space_4_sc_req(1 downto 1),
      memory_space_4_sc_ack => memory_space_4_sc_ack(1 downto 1),
      memory_space_4_sc_tag => memory_space_4_sc_tag(7 downto 4),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(6 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(6 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(31 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(21 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(7 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(20 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(3 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(1 downto 1),
      memory_space_8_sr_ack => memory_space_8_sr_ack(1 downto 1),
      memory_space_8_sr_addr => memory_space_8_sr_addr(1 downto 1),
      memory_space_8_sr_data => memory_space_8_sr_data(15 downto 8),
      memory_space_8_sr_tag => memory_space_8_sr_tag(43 downto 22),
      memory_space_8_sc_req => memory_space_8_sc_req(1 downto 1),
      memory_space_8_sc_ack => memory_space_8_sc_ack(1 downto 1),
      memory_space_8_sc_tag => memory_space_8_sc_tag(9 downto 5),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(21 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(4 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(20 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(7 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(6 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(1 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(6 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(21 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(4 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(20 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(7 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(21 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(7 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(4 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(21 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(4 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(7 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(21 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(20 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(3 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(7 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(21 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(4 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 2,
      addr_width => 1,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 1,
      num_stores => 2,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 2,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 2,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 1,
      num_stores => 2,
      addr_width => 1,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
