-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_711_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 : boolean;
  signal type_cast_711_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1040_inst_ack_0 : boolean;
  signal type_cast_711_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_ack_0 : boolean;
  signal type_cast_711_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1031_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1046_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1040_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1067_inst_ack_1 : boolean;
  signal phi_stmt_904_ack_0 : boolean;
  signal ptr_deref_602_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_992_inst_ack_1 : boolean;
  signal type_cast_594_inst_req_0 : boolean;
  signal addr_of_673_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_req_0 : boolean;
  signal WPIPE_Block1_start_992_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_req_1 : boolean;
  signal type_cast_558_inst_req_1 : boolean;
  signal array_obj_ref_672_index_offset_ack_1 : boolean;
  signal type_cast_558_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_518_inst_req_0 : boolean;
  signal type_cast_504_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_572_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_0 : boolean;
  signal ptr_deref_602_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 : boolean;
  signal array_obj_ref_672_index_offset_req_1 : boolean;
  signal type_cast_39_inst_req_0 : boolean;
  signal type_cast_39_inst_ack_0 : boolean;
  signal type_cast_39_inst_req_1 : boolean;
  signal type_cast_39_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 : boolean;
  signal type_cast_693_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_req_1 : boolean;
  signal WPIPE_Block0_start_980_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_0 : boolean;
  signal type_cast_52_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_1 : boolean;
  signal type_cast_52_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 : boolean;
  signal type_cast_558_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 : boolean;
  signal type_cast_693_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1028_inst_ack_0 : boolean;
  signal type_cast_680_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_req_0 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1049_inst_req_1 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal type_cast_558_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1049_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 : boolean;
  signal type_cast_1179_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 : boolean;
  signal type_cast_693_inst_req_1 : boolean;
  signal type_cast_680_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1046_inst_req_1 : boolean;
  signal type_cast_77_inst_req_0 : boolean;
  signal type_cast_77_inst_ack_0 : boolean;
  signal type_cast_77_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1040_inst_req_1 : boolean;
  signal type_cast_77_inst_ack_1 : boolean;
  signal addr_of_673_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 : boolean;
  signal addr_of_673_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 : boolean;
  signal type_cast_680_inst_ack_0 : boolean;
  signal array_obj_ref_672_index_offset_ack_0 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_1 : boolean;
  signal type_cast_89_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1040_inst_ack_1 : boolean;
  signal type_cast_89_inst_ack_0 : boolean;
  signal type_cast_89_inst_req_1 : boolean;
  signal type_cast_89_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1061_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 : boolean;
  signal type_cast_680_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_1 : boolean;
  signal type_cast_102_inst_req_0 : boolean;
  signal type_cast_102_inst_ack_0 : boolean;
  signal type_cast_102_inst_req_1 : boolean;
  signal type_cast_102_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1028_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1058_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_980_inst_req_0 : boolean;
  signal if_stmt_616_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 : boolean;
  signal array_obj_ref_672_index_offset_req_0 : boolean;
  signal WPIPE_Block0_start_980_inst_ack_0 : boolean;
  signal type_cast_114_inst_req_0 : boolean;
  signal type_cast_114_inst_ack_0 : boolean;
  signal type_cast_114_inst_req_1 : boolean;
  signal type_cast_114_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1052_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_req_1 : boolean;
  signal addr_of_673_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_1 : boolean;
  signal type_cast_127_inst_req_0 : boolean;
  signal type_cast_127_inst_ack_0 : boolean;
  signal type_cast_127_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_0 : boolean;
  signal type_cast_127_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1064_inst_req_1 : boolean;
  signal if_stmt_616_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal type_cast_317_inst_req_0 : boolean;
  signal type_cast_317_inst_ack_0 : boolean;
  signal type_cast_317_inst_req_1 : boolean;
  signal type_cast_317_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1061_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1055_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_326_inst_ack_1 : boolean;
  signal type_cast_1179_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_689_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_554_inst_req_0 : boolean;
  signal WPIPE_Block0_start_986_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1064_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_ack_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal type_cast_152_inst_req_0 : boolean;
  signal type_cast_152_inst_ack_0 : boolean;
  signal type_cast_152_inst_req_1 : boolean;
  signal WPIPE_Block0_start_980_inst_ack_1 : boolean;
  signal type_cast_152_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_707_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_992_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 : boolean;
  signal type_cast_693_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1046_inst_ack_1 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1046_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_req_1 : boolean;
  signal type_cast_177_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1001_inst_req_1 : boolean;
  signal type_cast_177_inst_ack_0 : boolean;
  signal type_cast_177_inst_req_1 : boolean;
  signal type_cast_177_inst_ack_1 : boolean;
  signal type_cast_540_inst_ack_1 : boolean;
  signal type_cast_540_inst_req_1 : boolean;
  signal if_stmt_616_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_0 : boolean;
  signal type_cast_189_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_1 : boolean;
  signal type_cast_189_inst_ack_1 : boolean;
  signal type_cast_540_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 : boolean;
  signal type_cast_540_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_590_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1028_inst_req_1 : boolean;
  signal type_cast_202_inst_req_0 : boolean;
  signal type_cast_202_inst_ack_0 : boolean;
  signal type_cast_202_inst_req_1 : boolean;
  signal type_cast_202_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1001_inst_req_0 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_504_inst_req_1 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1001_inst_ack_0 : boolean;
  signal type_cast_215_inst_req_0 : boolean;
  signal type_cast_215_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1061_inst_req_1 : boolean;
  signal type_cast_215_inst_req_1 : boolean;
  signal type_cast_215_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_986_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1028_inst_ack_1 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_req_1 : boolean;
  signal ptr_deref_602_store_0_ack_1 : boolean;
  signal type_cast_233_inst_req_0 : boolean;
  signal type_cast_233_inst_ack_0 : boolean;
  signal type_cast_233_inst_req_1 : boolean;
  signal type_cast_233_inst_ack_1 : boolean;
  signal ptr_deref_602_store_0_req_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal type_cast_237_inst_req_0 : boolean;
  signal type_cast_237_inst_ack_0 : boolean;
  signal type_cast_504_inst_ack_0 : boolean;
  signal type_cast_237_inst_req_1 : boolean;
  signal type_cast_237_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_536_inst_req_0 : boolean;
  signal type_cast_576_inst_ack_1 : boolean;
  signal type_cast_576_inst_req_1 : boolean;
  signal type_cast_241_inst_req_0 : boolean;
  signal type_cast_241_inst_ack_0 : boolean;
  signal type_cast_504_inst_req_0 : boolean;
  signal type_cast_241_inst_req_1 : boolean;
  signal type_cast_241_inst_ack_1 : boolean;
  signal type_cast_245_inst_req_0 : boolean;
  signal type_cast_245_inst_ack_0 : boolean;
  signal type_cast_245_inst_req_1 : boolean;
  signal type_cast_245_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1055_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_676_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal type_cast_576_inst_ack_0 : boolean;
  signal type_cast_576_inst_req_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal type_cast_522_inst_ack_1 : boolean;
  signal type_cast_522_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_req_1 : boolean;
  signal type_cast_594_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_276_inst_ack_1 : boolean;
  signal type_cast_280_inst_req_0 : boolean;
  signal type_cast_280_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1055_inst_req_1 : boolean;
  signal type_cast_280_inst_req_1 : boolean;
  signal type_cast_594_inst_req_1 : boolean;
  signal type_cast_280_inst_ack_1 : boolean;
  signal type_cast_522_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_ack_0 : boolean;
  signal type_cast_522_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_288_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_1 : boolean;
  signal WPIPE_Block0_start_983_inst_req_0 : boolean;
  signal type_cast_292_inst_req_0 : boolean;
  signal type_cast_292_inst_ack_0 : boolean;
  signal type_cast_292_inst_req_1 : boolean;
  signal type_cast_292_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_req_1 : boolean;
  signal type_cast_594_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_301_inst_ack_1 : boolean;
  signal type_cast_305_inst_req_0 : boolean;
  signal type_cast_305_inst_ack_0 : boolean;
  signal type_cast_305_inst_req_1 : boolean;
  signal type_cast_305_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_995_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_313_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_995_inst_ack_0 : boolean;
  signal type_cast_330_inst_req_0 : boolean;
  signal type_cast_330_inst_ack_0 : boolean;
  signal type_cast_330_inst_req_1 : boolean;
  signal type_cast_330_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_995_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1001_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_338_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_995_inst_ack_1 : boolean;
  signal type_cast_342_inst_req_0 : boolean;
  signal type_cast_342_inst_ack_0 : boolean;
  signal type_cast_342_inst_req_1 : boolean;
  signal type_cast_342_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_351_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal type_cast_355_inst_req_0 : boolean;
  signal type_cast_355_inst_ack_0 : boolean;
  signal type_cast_355_inst_req_1 : boolean;
  signal type_cast_355_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_998_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1043_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_363_inst_ack_1 : boolean;
  signal type_cast_367_inst_req_0 : boolean;
  signal type_cast_367_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_986_inst_req_1 : boolean;
  signal type_cast_367_inst_req_1 : boolean;
  signal type_cast_367_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1031_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1043_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_376_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_998_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal type_cast_380_inst_req_0 : boolean;
  signal type_cast_380_inst_ack_0 : boolean;
  signal type_cast_380_inst_req_1 : boolean;
  signal type_cast_380_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_998_inst_req_1 : boolean;
  signal WPIPE_Block0_start_986_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_998_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1052_inst_req_1 : boolean;
  signal if_stmt_394_branch_req_0 : boolean;
  signal if_stmt_394_branch_ack_1 : boolean;
  signal if_stmt_394_branch_ack_0 : boolean;
  signal if_stmt_409_branch_req_0 : boolean;
  signal if_stmt_409_branch_ack_1 : boolean;
  signal if_stmt_409_branch_ack_0 : boolean;
  signal type_cast_436_inst_req_0 : boolean;
  signal type_cast_436_inst_ack_0 : boolean;
  signal type_cast_436_inst_req_1 : boolean;
  signal type_cast_436_inst_ack_1 : boolean;
  signal array_obj_ref_465_index_offset_req_0 : boolean;
  signal array_obj_ref_465_index_offset_ack_0 : boolean;
  signal array_obj_ref_465_index_offset_req_1 : boolean;
  signal array_obj_ref_465_index_offset_ack_1 : boolean;
  signal addr_of_466_final_reg_req_0 : boolean;
  signal addr_of_466_final_reg_ack_0 : boolean;
  signal addr_of_466_final_reg_req_1 : boolean;
  signal addr_of_466_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_469_inst_ack_1 : boolean;
  signal type_cast_473_inst_req_0 : boolean;
  signal type_cast_473_inst_ack_0 : boolean;
  signal type_cast_473_inst_req_1 : boolean;
  signal type_cast_473_inst_ack_1 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_482_inst_ack_1 : boolean;
  signal type_cast_486_inst_req_0 : boolean;
  signal type_cast_486_inst_ack_0 : boolean;
  signal type_cast_486_inst_req_1 : boolean;
  signal type_cast_486_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_500_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_725_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1058_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1055_inst_req_0 : boolean;
  signal type_cast_729_inst_req_0 : boolean;
  signal type_cast_729_inst_ack_0 : boolean;
  signal type_cast_729_inst_req_1 : boolean;
  signal type_cast_729_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1061_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1067_inst_req_1 : boolean;
  signal WPIPE_Block1_start_992_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1049_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_743_inst_ack_1 : boolean;
  signal type_cast_1247_inst_ack_1 : boolean;
  signal type_cast_747_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1037_inst_ack_1 : boolean;
  signal type_cast_747_inst_ack_0 : boolean;
  signal type_cast_747_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1037_inst_req_1 : boolean;
  signal type_cast_747_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1049_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_761_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1058_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1058_inst_req_0 : boolean;
  signal type_cast_765_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1037_inst_ack_0 : boolean;
  signal type_cast_765_inst_ack_0 : boolean;
  signal type_cast_765_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1037_inst_req_0 : boolean;
  signal type_cast_765_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1010_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_779_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1010_inst_req_1 : boolean;
  signal type_cast_783_inst_req_0 : boolean;
  signal type_cast_783_inst_ack_0 : boolean;
  signal type_cast_783_inst_req_1 : boolean;
  signal type_cast_783_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1067_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1010_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_989_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_797_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_989_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1064_inst_ack_0 : boolean;
  signal if_stmt_1304_branch_ack_1 : boolean;
  signal type_cast_801_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1034_inst_ack_1 : boolean;
  signal type_cast_801_inst_ack_0 : boolean;
  signal type_cast_801_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1034_inst_req_1 : boolean;
  signal type_cast_801_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1067_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_0 : boolean;
  signal phi_stmt_904_req_0 : boolean;
  signal WPIPE_Block3_start_1064_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1034_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1034_inst_req_0 : boolean;
  signal ptr_deref_809_store_0_req_0 : boolean;
  signal ptr_deref_809_store_0_ack_0 : boolean;
  signal ptr_deref_809_store_0_req_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_ack_1 : boolean;
  signal ptr_deref_809_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1052_inst_req_0 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_1 : boolean;
  signal if_stmt_823_branch_req_0 : boolean;
  signal WPIPE_Block0_start_983_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1025_inst_ack_1 : boolean;
  signal if_stmt_823_branch_ack_1 : boolean;
  signal WPIPE_Block2_start_1025_inst_req_1 : boolean;
  signal if_stmt_823_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1007_inst_ack_0 : boolean;
  signal type_cast_834_inst_req_0 : boolean;
  signal type_cast_834_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1025_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_983_inst_ack_0 : boolean;
  signal type_cast_834_inst_req_1 : boolean;
  signal type_cast_834_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1043_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1007_inst_req_0 : boolean;
  signal type_cast_838_inst_req_0 : boolean;
  signal type_cast_838_inst_ack_0 : boolean;
  signal type_cast_838_inst_req_1 : boolean;
  signal type_cast_838_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_989_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_989_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1043_inst_req_1 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal type_cast_1267_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1025_inst_req_0 : boolean;
  signal if_stmt_860_branch_req_0 : boolean;
  signal if_stmt_860_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_977_inst_ack_1 : boolean;
  signal if_stmt_860_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1031_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1004_inst_ack_1 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1031_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_977_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1052_inst_ack_1 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1004_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1004_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1004_inst_req_0 : boolean;
  signal array_obj_ref_916_index_offset_req_0 : boolean;
  signal array_obj_ref_916_index_offset_ack_0 : boolean;
  signal array_obj_ref_916_index_offset_req_1 : boolean;
  signal array_obj_ref_916_index_offset_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 : boolean;
  signal addr_of_917_final_reg_req_0 : boolean;
  signal addr_of_917_final_reg_ack_0 : boolean;
  signal addr_of_917_final_reg_req_1 : boolean;
  signal addr_of_917_final_reg_ack_1 : boolean;
  signal if_stmt_1304_branch_ack_0 : boolean;
  signal type_cast_1257_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 : boolean;
  signal type_cast_1257_inst_ack_0 : boolean;
  signal ptr_deref_920_store_0_req_0 : boolean;
  signal ptr_deref_920_store_0_ack_0 : boolean;
  signal ptr_deref_920_store_0_req_1 : boolean;
  signal ptr_deref_920_store_0_ack_1 : boolean;
  signal type_cast_1267_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1272_inst_ack_1 : boolean;
  signal if_stmt_935_branch_req_0 : boolean;
  signal type_cast_1267_inst_ack_1 : boolean;
  signal if_stmt_935_branch_ack_1 : boolean;
  signal if_stmt_935_branch_ack_0 : boolean;
  signal call_stmt_946_call_req_0 : boolean;
  signal call_stmt_946_call_ack_0 : boolean;
  signal call_stmt_946_call_req_1 : boolean;
  signal call_stmt_946_call_ack_1 : boolean;
  signal type_cast_1179_inst_req_1 : boolean;
  signal type_cast_951_inst_req_0 : boolean;
  signal type_cast_951_inst_ack_0 : boolean;
  signal type_cast_951_inst_req_1 : boolean;
  signal type_cast_951_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_953_inst_req_0 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_953_inst_req_1 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_956_inst_req_0 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_956_inst_req_1 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_959_inst_req_0 : boolean;
  signal WPIPE_Block0_start_959_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_959_inst_req_1 : boolean;
  signal WPIPE_Block0_start_959_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_962_inst_req_0 : boolean;
  signal WPIPE_Block0_start_962_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_962_inst_req_1 : boolean;
  signal WPIPE_Block0_start_962_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_965_inst_req_0 : boolean;
  signal WPIPE_Block0_start_965_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_965_inst_req_1 : boolean;
  signal WPIPE_Block0_start_965_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_968_inst_req_0 : boolean;
  signal WPIPE_Block0_start_968_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_968_inst_req_1 : boolean;
  signal WPIPE_Block0_start_968_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_971_inst_req_0 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_971_inst_req_1 : boolean;
  signal WPIPE_Block0_start_971_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_974_inst_req_0 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_974_inst_req_1 : boolean;
  signal WPIPE_Block0_start_974_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_977_inst_req_0 : boolean;
  signal WPIPE_Block0_start_977_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1070_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1070_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1070_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1070_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1073_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1073_inst_ack_0 : boolean;
  signal type_cast_1267_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1073_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1073_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1284_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_req_0 : boolean;
  signal phi_stmt_453_ack_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1076_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1076_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1079_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1079_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1079_inst_req_1 : boolean;
  signal phi_stmt_453_req_1 : boolean;
  signal WPIPE_Block3_start_1079_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1082_inst_req_0 : boolean;
  signal type_cast_459_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1082_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1082_inst_req_1 : boolean;
  signal type_cast_459_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1082_inst_ack_1 : boolean;
  signal phi_stmt_904_req_1 : boolean;
  signal WPIPE_Block3_start_1085_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1085_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1085_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1085_inst_ack_1 : boolean;
  signal type_cast_910_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1088_inst_req_0 : boolean;
  signal type_cast_459_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1088_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1088_inst_req_1 : boolean;
  signal type_cast_459_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1088_inst_ack_1 : boolean;
  signal type_cast_910_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1091_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1091_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1091_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1091_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1094_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1094_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1094_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1094_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1098_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1098_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1098_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1098_inst_ack_1 : boolean;
  signal type_cast_910_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1101_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1101_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1269_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1101_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1101_inst_ack_1 : boolean;
  signal phi_stmt_1176_ack_0 : boolean;
  signal type_cast_910_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1104_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1104_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1104_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1104_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1107_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1107_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1107_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1281_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1107_inst_ack_1 : boolean;
  signal call_stmt_1111_call_req_0 : boolean;
  signal call_stmt_1111_call_ack_0 : boolean;
  signal type_cast_1179_inst_req_0 : boolean;
  signal call_stmt_1111_call_req_1 : boolean;
  signal phi_stmt_453_req_0 : boolean;
  signal call_stmt_1111_call_ack_1 : boolean;
  signal type_cast_1247_inst_req_1 : boolean;
  signal type_cast_1115_inst_req_0 : boolean;
  signal type_cast_1115_inst_ack_0 : boolean;
  signal if_stmt_1304_branch_req_0 : boolean;
  signal type_cast_1115_inst_req_1 : boolean;
  signal type_cast_1115_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1122_inst_ack_1 : boolean;
  signal if_stmt_1132_branch_req_0 : boolean;
  signal if_stmt_1132_branch_ack_1 : boolean;
  signal if_stmt_1132_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_ack_0 : boolean;
  signal type_cast_1159_inst_req_0 : boolean;
  signal type_cast_1159_inst_ack_0 : boolean;
  signal type_cast_1159_inst_req_1 : boolean;
  signal type_cast_1159_inst_ack_1 : boolean;
  signal phi_stmt_1176_req_0 : boolean;
  signal phi_stmt_660_ack_0 : boolean;
  signal phi_stmt_660_req_0 : boolean;
  signal type_cast_1257_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_ack_1 : boolean;
  signal array_obj_ref_1188_index_offset_req_0 : boolean;
  signal array_obj_ref_1188_index_offset_ack_0 : boolean;
  signal array_obj_ref_1188_index_offset_req_1 : boolean;
  signal array_obj_ref_1188_index_offset_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_req_1 : boolean;
  signal addr_of_1189_final_reg_req_0 : boolean;
  signal addr_of_1189_final_reg_ack_0 : boolean;
  signal addr_of_1189_final_reg_req_1 : boolean;
  signal addr_of_1189_final_reg_ack_1 : boolean;
  signal type_cast_663_inst_ack_1 : boolean;
  signal type_cast_663_inst_req_1 : boolean;
  signal type_cast_663_inst_ack_0 : boolean;
  signal type_cast_663_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_req_0 : boolean;
  signal ptr_deref_1193_load_0_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1278_inst_req_0 : boolean;
  signal ptr_deref_1193_load_0_ack_0 : boolean;
  signal type_cast_1257_inst_req_1 : boolean;
  signal ptr_deref_1193_load_0_req_1 : boolean;
  signal ptr_deref_1193_load_0_ack_1 : boolean;
  signal type_cast_1197_inst_req_0 : boolean;
  signal type_cast_1197_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 : boolean;
  signal type_cast_1197_inst_req_1 : boolean;
  signal type_cast_1197_inst_ack_1 : boolean;
  signal type_cast_1247_inst_ack_0 : boolean;
  signal type_cast_1207_inst_req_0 : boolean;
  signal type_cast_1207_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_0 : boolean;
  signal phi_stmt_1176_req_1 : boolean;
  signal type_cast_1207_inst_req_1 : boolean;
  signal type_cast_1207_inst_ack_1 : boolean;
  signal type_cast_1247_inst_req_0 : boolean;
  signal type_cast_1217_inst_req_0 : boolean;
  signal type_cast_1217_inst_ack_0 : boolean;
  signal type_cast_1217_inst_req_1 : boolean;
  signal type_cast_1217_inst_ack_1 : boolean;
  signal type_cast_1227_inst_req_0 : boolean;
  signal type_cast_1227_inst_ack_0 : boolean;
  signal type_cast_1227_inst_req_1 : boolean;
  signal type_cast_1227_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1275_inst_ack_1 : boolean;
  signal phi_stmt_660_req_1 : boolean;
  signal type_cast_1237_inst_req_0 : boolean;
  signal type_cast_1237_inst_ack_0 : boolean;
  signal type_cast_1237_inst_req_1 : boolean;
  signal type_cast_1237_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(425 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(425);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_33/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/branch_block_stmt_33__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393__entry__
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_update_start_
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/cr
      -- 
    rr_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_0); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_39_inst_req_1); -- 
    cr_182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_52_inst_req_1); -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_64_inst_req_1); -- 
    cr_238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_77_inst_req_1); -- 
    cr_266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_89_inst_req_1); -- 
    cr_294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_102_inst_req_1); -- 
    cr_322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_114_inst_req_1); -- 
    cr_350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_127_inst_req_1); -- 
    cr_756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_317_inst_req_1); -- 
    cr_378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_139_inst_req_1); -- 
    cr_406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_152_inst_req_1); -- 
    cr_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_164_inst_req_1); -- 
    cr_462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_177_inst_req_1); -- 
    cr_490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_189_inst_req_1); -- 
    cr_518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_202_inst_req_1); -- 
    cr_532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_215_inst_req_1); -- 
    cr_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_219_inst_req_1); -- 
    cr_574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_233_inst_req_1); -- 
    cr_588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_237_inst_req_1); -- 
    cr_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_241_inst_req_1); -- 
    cr_616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_245_inst_req_1); -- 
    cr_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_267_inst_req_1); -- 
    cr_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_280_inst_req_1); -- 
    cr_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_292_inst_req_1); -- 
    cr_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_305_inst_req_1); -- 
    cr_784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_330_inst_req_1); -- 
    cr_812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_342_inst_req_1); -- 
    cr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_355_inst_req_1); -- 
    cr_868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_367_inst_req_1); -- 
    cr_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_380_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_update_start_
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/cr
      -- 
    ra_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_35_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_35_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/rr
      -- 
    ca_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_35_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_39_inst_req_0); -- 
    rr_163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Sample/ra
      -- 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_39_Update/ca
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_39_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_update_start_
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/cr
      -- 
    ra_164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_48_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_48_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/rr
      -- 
    ca_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_48_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_52_inst_req_0); -- 
    rr_191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Sample/ra
      -- 
    ra_178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_52_Update/ca
      -- 
    ca_183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_update_start_
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/cr
      -- 
    ra_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_60_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_60_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/rr
      -- 
    ca_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_60_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_64_inst_req_0); -- 
    rr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_64_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_update_start_
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/cr
      -- 
    ra_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_73_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_73_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/rr
      -- 
    ca_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_73_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_77_inst_req_0); -- 
    rr_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Sample/ra
      -- 
    ra_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_77_Update/ca
      -- 
    ca_239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_update_start_
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/cr
      -- 
    ra_248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_85_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_85_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/rr
      -- 
    ca_253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_85_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_89_inst_req_0); -- 
    rr_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Sample/ra
      -- 
    ra_262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_89_Update/ca
      -- 
    ca_267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_89_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_update_start_
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/cr
      -- 
    ra_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_98_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_98_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/rr
      -- 
    ca_281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_98_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_102_inst_req_0); -- 
    rr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Sample/ra
      -- 
    ra_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_102_Update/ca
      -- 
    ca_295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_102_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_update_start_
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/cr
      -- 
    ra_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_110_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_110_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/rr
      -- 
    ca_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_110_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_114_inst_req_0); -- 
    rr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Sample/ra
      -- 
    ra_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_114_Update/ca
      -- 
    ca_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_114_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_update_start_
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/cr
      -- 
    ra_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_123_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_sample_start_
      -- 
    ca_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_127_inst_req_0); -- 
    rr_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Sample/ra
      -- 
    ra_346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_127_Update/ca
      -- 
    ca_351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_update_start_
      -- 
    ra_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_135_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_135_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/rr
      -- 
    ca_365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_135_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_139_inst_req_0); -- 
    rr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Sample/ra
      -- 
    ra_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_139_Update/ca
      -- 
    ca_379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_update_start_
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/cr
      -- 
    ra_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_148_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_148_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/rr
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_148_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_0); -- 
    rr_401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_152_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Sample/ra
      -- 
    ra_402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_152_Update/ca
      -- 
    ca_407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_152_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_update_start_
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/cr
      -- 
    ra_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_160_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_160_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/rr
      -- 
    ca_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_160_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_164_inst_req_0); -- 
    rr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Sample/ra
      -- 
    ra_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_164_Update/ca
      -- 
    ca_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_update_start_
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/cr
      -- 
    ra_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_173_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_173_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/rr
      -- 
    ca_449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_173_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_177_inst_req_0); -- 
    rr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Sample/ra
      -- 
    ra_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_177_Update/ca
      -- 
    ca_463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_177_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_update_start_
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/cr
      -- 
    ra_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_185_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_185_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/rr
      -- 
    ca_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_185_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_0); -- 
    rr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_189_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Sample/ra
      -- 
    ra_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_189_Update/ca
      -- 
    ca_491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_update_start_
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/cr
      -- 
    ra_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_198_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_198_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/rr
      -- 
    ca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_198_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_202_inst_req_0); -- 
    rr_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_263_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Sample/ra
      -- 
    ra_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_202_Update/ca
      -- 
    ca_519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_202_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/rr
      -- 
    rr_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_211_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Sample/ra
      -- 
    ra_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_211_Update/ca
      -- 
    ca_533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/rr
      -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_215_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Sample/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_215_Update/ca
      -- 
    ca_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_215_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/rr
      -- 
    rr_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_219_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Sample/ra
      -- 
    ra_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_219_Update/ca
      -- 
    ca_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/rr
      -- 
    rr_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_233_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Sample/ra
      -- 
    ra_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_233_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_233_Update/ca
      -- 
    ca_575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_233_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/rr
      -- 
    rr_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_237_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Sample/ra
      -- 
    ra_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_237_Update/ca
      -- 
    ca_589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: 	44 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/rr
      -- 
    rr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_241_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(48) & convTranspose_CP_39_elements(44);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Sample/ra
      -- 
    ra_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_241_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_241_Update/ca
      -- 
    ca_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_241_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/rr
      -- 
    rr_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_245_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Sample/ra
      -- 
    ra_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_245_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_245_Update/ca
      -- 
    ca_617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_245_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_update_start_
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/cr
      -- 
    ra_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_263_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_263_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_263_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/rr
      -- 
    ca_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_263_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_267_inst_req_0); -- 
    rr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_276_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Sample/ra
      -- 
    ra_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_267_Update/ca
      -- 
    ca_645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_update_start_
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/cr
      -- 
    ra_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_276_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_276_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_276_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/rr
      -- 
    ca_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_276_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_280_inst_req_0); -- 
    rr_681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_288_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Sample/ra
      -- 
    ra_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_280_Update/ca
      -- 
    ca_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_update_start_
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/cr
      -- 
    ra_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_288_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_288_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_288_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/rr
      -- 
    ca_687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_288_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_292_inst_req_0); -- 
    rr_709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_301_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Sample/ra
      -- 
    ra_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_292_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_292_Update/ca
      -- 
    ca_701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_292_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_update_start_
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/cr
      -- 
    ra_710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_301_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_301_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_301_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/rr
      -- 
    ca_715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_301_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_305_inst_req_0); -- 
    rr_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_313_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Sample/ra
      -- 
    ra_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_305_Update/ca
      -- 
    ca_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_update_start_
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/cr
      -- 
    ra_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_313_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_313_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_313_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_sample_start_
      -- 
    ca_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_313_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_317_inst_req_0); -- 
    rr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_326_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_sample_completed_
      -- 
    ra_752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_317_Update/ca
      -- 
    ca_757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_317_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_update_start_
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/cr
      -- 
    ra_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_326_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_326_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_326_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/rr
      -- 
    ca_771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_326_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_330_inst_req_0); -- 
    rr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_338_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Sample/ra
      -- 
    ra_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_330_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_330_Update/ca
      -- 
    ca_785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_330_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_update_start_
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/cr
      -- 
    ra_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_338_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_338_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_338_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/rr
      -- 
    ca_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_338_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_342_inst_req_0); -- 
    rr_821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_351_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Sample/ra
      -- 
    ra_808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_342_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_342_Update/ca
      -- 
    ca_813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_342_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_update_start_
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/cr
      -- 
    ra_822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_351_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_351_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_351_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/rr
      -- 
    ca_827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_351_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_355_inst_req_0); -- 
    rr_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_363_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Sample/ra
      -- 
    ra_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_355_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_355_Update/ca
      -- 
    ca_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_355_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_update_start_
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/cr
      -- 
    ra_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_363_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_363_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_363_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/rr
      -- 
    ca_855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_363_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_367_inst_req_0); -- 
    rr_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_376_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Sample/ra
      -- 
    ra_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_367_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_367_Update/ca
      -- 
    ca_869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_367_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_update_start_
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/cr
      -- 
    ra_878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_376_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_376_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/RPIPE_ConvTranspose_input_pipe_376_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/rr
      -- 
    ca_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_376_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_380_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Sample/ra
      -- 
    ra_892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/type_cast_380_Update/ca
      -- 
    ca_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393__exit__
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394__entry__
      -- CP-element group 118: 	 branch_block_stmt_33/assign_stmt_36_to_assign_stmt_393/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_33/R_cmp417_395_place
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_33/if_stmt_394_else_link/$entry
      -- 
    branch_req_905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_394_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415__exit__
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450__entry__
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_394_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/if_stmt_394_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph419
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_update_start_
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiAck/dummy
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/merge_stmt_415_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph419_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_33/entry_bbx_xnph419_PhiReq/$entry
      -- 
    if_choice_transition_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_394_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_436_inst_req_0); -- 
    cr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_436_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	398 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_394_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/if_stmt_394_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond176x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond176x_xpreheader_PhiReq/$exit
      -- CP-element group 120: 	 branch_block_stmt_33/entry_forx_xcond176x_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_394_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	398 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622__exit__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657__entry__
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_update_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiAck/dummy
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_bbx_xnph415_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_bbx_xnph415_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_409_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_33/if_stmt_409_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_bbx_xnph415
      -- CP-element group 121: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_33/merge_stmt_622_PhiReqMerge
      -- 
    if_choice_transition_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_409_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    rr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_643_inst_req_0); -- 
    cr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_643_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	398 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	411 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_409_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/if_stmt_409_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_forx_xend236
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_forx_xend236_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_33/forx_xcond176x_xpreheader_forx_xend236_PhiReq/$entry
      -- 
    else_choice_transition_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_409_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Sample/ra
      -- 
    ra_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	399 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450__exit__
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_33/assign_stmt_421_to_assign_stmt_450/type_cast_436_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/$entry
      -- CP-element group 124: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/$entry
      -- 
    ca_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	404 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/ack
      -- 
    ack_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_465_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	404 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/req
      -- 
    ack_989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_465_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_466_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_request/ack
      -- 
    ack_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_466_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	404 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/ack
      -- 
    ack_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_466_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	404 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_update_start_
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/cr
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_469_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_469_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/rr
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_469_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_473_inst_req_0); -- 
    rr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_482_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Sample/ra
      -- 
    ra_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	404 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/ca
      -- 
    ca_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_update_start_
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/cr
      -- 
    ra_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_482_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_482_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_482_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/rr
      -- 
    ca_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_482_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_486_inst_req_0); -- 
    rr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_500_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Sample/ra
      -- 
    ra_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	404 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/ca
      -- 
    ca_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_update_start_
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/cr
      -- 
    ra_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_500_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_500_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_500_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/$entry
      -- 
    ca_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_500_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_504_inst_req_0); -- 
    rr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_518_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_sample_completed_
      -- 
    ra_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	404 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_update_completed_
      -- 
    ca_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_update_start_
      -- CP-element group 141: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_sample_completed_
      -- 
    ra_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_518_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_518_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_518_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/$entry
      -- 
    ca_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_518_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_522_inst_req_0); -- 
    rr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_536_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Sample/$exit
      -- 
    ra_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_522_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	404 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_update_completed_
      -- 
    ca_1116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_522_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_update_start_
      -- CP-element group 145: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_sample_completed_
      -- 
    ra_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_536_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_536_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_536_update_completed_
      -- 
    ca_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_536_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_540_inst_req_0); -- 
    rr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_554_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_sample_completed_
      -- 
    ra_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	404 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_update_completed_
      -- 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_update_start_
      -- CP-element group 149: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_sample_completed_
      -- 
    ra_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_554_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_554_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_554_update_completed_
      -- 
    ca_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_554_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_558_inst_req_0); -- 
    rr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_572_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_sample_completed_
      -- 
    ra_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_558_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	404 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_update_completed_
      -- 
    ca_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_558_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_update_start_
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Sample/$exit
      -- 
    ra_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_572_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_572_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_572_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/$entry
      -- 
    ca_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_572_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_576_inst_req_0); -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_590_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Sample/$exit
      -- 
    ra_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_576_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	404 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_update_completed_
      -- 
    ca_1200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_576_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_update_start_
      -- CP-element group 157: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_sample_completed_
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_590_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_590_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_590_update_completed_
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_590_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_594_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Sample/ra
      -- 
    ra_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_594_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	404 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/$exit
      -- 
    ca_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_594_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/ptr_deref_602_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_sample_start_
      -- 
    rr_1266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_602_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(156);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_sample_completed_
      -- 
    ra_1267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	404 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/$exit
      -- 
    ca_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615__exit__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616__entry__
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/R_exitcond3_617_place
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/if_stmt_616_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/$exit
      -- 
    branch_req_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_616_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	398 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400__exit__
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_616_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_33/if_stmt_616_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xcond176x_xpreheaderx_xloopexit_forx_xcond176x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/merge_stmt_400_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_33/forx_xbody_forx_xcond176x_xpreheaderx_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_616_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	400 
    -- CP-element group 166: 	401 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_616_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_33/if_stmt_616_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/cr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/$entry
      -- CP-element group 166: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_1295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_616_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    cr_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_459_inst_req_1); -- 
    rr_3105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_459_inst_req_0); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Sample/$exit
      -- 
    ra_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	405 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657__exit__
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/$exit
      -- CP-element group 168: 	 branch_block_stmt_33/assign_stmt_628_to_assign_stmt_657/type_cast_643_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/$entry
      -- CP-element group 168: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$entry
      -- 
    ca_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	410 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_sample_complete
      -- 
    ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	410 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_sample_start_
      -- 
    ack_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_673_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_request/ack
      -- CP-element group 171: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_sample_completed_
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_673_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	410 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_word_addrgen/root_register_ack
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_673_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	410 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_update_start_
      -- CP-element group 173: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_sample_completed_
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_676_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_676_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	177 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_update_completed_
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_676_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_680_inst_req_0); -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_689_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Sample/$exit
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	410 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_update_completed_
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_update_start_
      -- CP-element group 177: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_sample_completed_
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_689_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_689_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_689_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/$entry
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_689_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_693_inst_req_0); -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_707_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Sample/$exit
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	410 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_update_completed_
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_update_start_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Sample/ra
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_707_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_707_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_707_Update/$exit
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_707_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_711_inst_req_0); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_725_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Sample/$exit
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_711_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	410 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/$exit
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_711_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_update_start_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/cr
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_725_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_725_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_725_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/rr
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_725_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_729_inst_req_0); -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_743_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Sample/ra
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_729_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	410 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/ca
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_729_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_update_start_
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/cr
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_743_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_743_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_743_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/rr
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_743_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_747_inst_req_0); -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_761_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Sample/ra
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	410 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/ca
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_747_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_update_start_
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/cr
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_761_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_761_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_761_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/rr
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_761_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_765_inst_req_0); -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_779_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Sample/ra
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_765_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	410 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_765_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_update_start_
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/cr
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_779_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_779_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_779_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/rr
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_779_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_783_inst_req_0); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_797_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Sample/ra
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	410 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/ca
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_update_start_
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/cr
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_797_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_797_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_797_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/rr
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_797_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_801_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Sample/ra
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	410 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/ca
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/ptr_deref_809_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/rr
      -- 
    rr_1625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_809_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204) & convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Sample/word_access_start/word_0/ra
      -- 
    ra_1626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_809_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	410 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/ca
      -- 
    ca_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_809_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822__exit__
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823__entry__
      -- CP-element group 208: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_33/R_exitcond2_824_place
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_33/if_stmt_823_else_link/$entry
      -- 
    branch_req_1645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_823_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(207) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	411 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829__exit__
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend236x_xloopexit_forx_xend236
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_823_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/if_stmt_823_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody182_forx_xend236x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend236x_xloopexit_forx_xend236_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xend236x_xloopexit_forx_xend236_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/merge_stmt_829_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody182_forx_xend236x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_33/forx_xbody182_forx_xend236x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_823_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	406 
    -- CP-element group 210: 	407 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_823_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_33/if_stmt_823_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/$entry
      -- CP-element group 210: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/$entry
      -- 
    else_choice_transition_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_823_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    cr_3164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_663_inst_req_1); -- 
    rr_3159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_663_inst_req_0); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	411 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/ra
      -- 
    ra_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_834_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	411 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/ca
      -- 
    ca_1673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_834_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	411 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/ra
      -- 
    ra_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	411 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/ca
      -- 
    ca_1687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	411 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/ra
      -- 
    ra_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	411 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/ca
      -- 
    ca_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859__exit__
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860__entry__
      -- CP-element group 217: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_33/R_cmp250409_861_place
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_33/if_stmt_860_else_link/$entry
      -- 
    branch_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_860_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866__exit__
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901__entry__
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_860_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/if_stmt_860_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend236_bbx_xnph411
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_update_start_
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/merge_stmt_866_PhiAck/dummy
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend236_bbx_xnph411_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_33/forx_xend236_bbx_xnph411_PhiReq/$entry
      -- 
    if_choice_transition_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_860_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_887_inst_req_0); -- 
    cr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_887_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	418 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend236_forx_xend259_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend236_forx_xend259_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_860_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_33/if_stmt_860_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_33/forx_xend236_forx_xend259
      -- 
    else_choice_transition_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_860_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Sample/ra
      -- 
    ra_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	412 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901__exit__
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_33/assign_stmt_872_to_assign_stmt_901/type_cast_887_Update/ca
      -- 
    ca_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	417 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/ack
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_916_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	417 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/req
      -- 
    ack_1771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_916_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_917_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_request/ack
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_917_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	417 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/ptr_deref_920_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/rr
      -- 
    ack_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_917_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_920_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Sample/word_access_start/word_0/ra
      -- 
    ra_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_920_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	417 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/ca
      -- 
    ca_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_920_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934__exit__
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935__entry__
      -- CP-element group 228: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_33/R_exitcond_936_place
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_33/if_stmt_935_else_link/$entry
      -- 
    branch_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_935_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	418 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941__exit__
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend259x_xloopexit_forx_xend259
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend259x_xloopexit_forx_xend259_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/merge_stmt_941_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody252_forx_xend259x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody252_forx_xend259x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_935_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_33/if_stmt_935_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xbody252_forx_xend259x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_33/forx_xend259x_xloopexit_forx_xend259_PhiReq/$entry
      -- 
    if_choice_transition_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_935_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	413 
    -- CP-element group 230: 	414 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_935_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_33/if_stmt_935_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/cr
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/$entry
      -- 
    else_choice_transition_1853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_935_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    cr_3241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_910_inst_req_1); -- 
    rr_3236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_910_inst_req_0); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	418 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/cra
      -- 
    cra_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_946_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	418 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/rr
      -- 
    cca_1872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_946_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_951_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Sample/ra
      -- 
    ra_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_951_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	418 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	339 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/ca
      -- 
    ca_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_951_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	418 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_update_start_
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/req
      -- 
    ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_953_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/req
      -- 
    ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_956_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_update_start_
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/req
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_956_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_956_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/req
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_959_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_update_start_
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/req
      -- 
    ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_959_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_959_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_959_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/req
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_959_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_962_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_update_start_
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/req
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_962_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_962_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_962_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/req
      -- 
    ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_962_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_965_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_update_start_
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/req
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_965_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_965_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_965_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/req
      -- 
    ack_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_965_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_968_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_update_start_
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/req
      -- 
    ack_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_968_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_968_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_968_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/req
      -- 
    ack_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_968_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_971_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_update_start_
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/req
      -- 
    ack_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_971_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_971_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/req
      -- 
    ack_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_971_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_974_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_update_start_
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/req
      -- 
    ack_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_974_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_974_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/req
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_974_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_977_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/req
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_update_start_
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Sample/ack
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_977_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_977_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_977_update_completed_
      -- 
    ack_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_977_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_980_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/req
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_update_start_
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_sample_completed_
      -- 
    ack_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_980_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_980_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_980_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/req
      -- 
    ack_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_980_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_983_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_update_start_
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/req
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Sample/ack
      -- 
    ack_2035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_983_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_983_Update/$exit
      -- 
    ack_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_983_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_986_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_update_start_
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/req
      -- 
    ack_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_986_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_986_inst_req_1); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	339 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_986_Update/ack
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_986_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	418 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/req
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_update_start_
      -- CP-element group 259: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_sample_completed_
      -- 
    ack_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_989_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block1_start_989_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_update_completed_
      -- 
    ack_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_989_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block1_start_992_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/req
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_update_start_
      -- CP-element group 261: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_sample_completed_
      -- 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_992_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block1_start_992_inst_req_1); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/req
      -- CP-element group 262: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_992_update_completed_
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_992_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    req_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(262), ack => WPIPE_Block1_start_995_inst_req_0); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_update_start_
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/req
      -- 
    ack_2091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_995_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_995_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_995_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/req
      -- 
    ack_2096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_995_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_998_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_update_start_
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/req
      -- 
    ack_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_998_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_998_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_998_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/$entry
      -- 
    ack_2110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_998_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1001_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/req
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_update_start_
      -- CP-element group 267: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_sample_completed_
      -- 
    ack_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1001_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1001_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1001_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/$entry
      -- 
    ack_2124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1001_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1004_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/req
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_update_start_
      -- 
    ack_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1004_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1004_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1004_update_completed_
      -- 
    ack_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1004_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1007_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/req
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_update_start_
      -- CP-element group 271: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_sample_completed_
      -- 
    ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1007_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1007_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1007_update_completed_
      -- 
    ack_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1007_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1010_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/req
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_update_start_
      -- CP-element group 273: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_sample_completed_
      -- 
    ack_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1010_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1010_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1010_update_completed_
      -- 
    ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1010_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1013_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/req
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_update_start_
      -- CP-element group 275: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_sample_completed_
      -- 
    ack_2175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1013_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1013_update_completed_
      -- 
    ack_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1016_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/req
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_update_start_
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_sample_completed_
      -- 
    ack_2189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1016_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1016_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/req
      -- 
    ack_2194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_update_start_
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/req
      -- 
    ack_2203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 280:  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/req
      -- 
    ack_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    req_2216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(280), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/req
      -- 
    ack_2217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    req_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(281), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	339 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_1022_Update/ack
      -- 
    ack_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	418 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_update_start_
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/req
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/ack
      -- CP-element group 283: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/$exit
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1025_inst_ack_0, ack => convTranspose_CP_39_elements(283)); -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block2_start_1025_inst_req_1); -- 
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/req
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_update_completed_
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1025_inst_ack_1, ack => convTranspose_CP_39_elements(284)); -- 
    req_2244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block2_start_1028_inst_req_0); -- 
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/req
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_update_start_
      -- CP-element group 285: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_sample_completed_
      -- 
    ack_2245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1028_inst_ack_0, ack => convTranspose_CP_39_elements(285)); -- 
    req_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(285), ack => WPIPE_Block2_start_1028_inst_req_1); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1028_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/req
      -- 
    ack_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1028_inst_ack_1, ack => convTranspose_CP_39_elements(286)); -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(286), ack => WPIPE_Block2_start_1031_inst_req_0); -- 
    -- CP-element group 287:  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_update_start_
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/req
      -- CP-element group 287: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/$entry
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1031_inst_ack_0, ack => convTranspose_CP_39_elements(287)); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(287), ack => WPIPE_Block2_start_1031_inst_req_1); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1031_Update/$exit
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1031_inst_ack_1, ack => convTranspose_CP_39_elements(288)); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block2_start_1034_inst_req_0); -- 
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/req
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_update_start_
      -- CP-element group 289: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_sample_completed_
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1034_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block2_start_1034_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1034_update_completed_
      -- 
    ack_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1034_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block2_start_1037_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/req
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_update_start_
      -- CP-element group 291: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_sample_completed_
      -- 
    ack_2287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1037_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block2_start_1037_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1037_update_completed_
      -- 
    ack_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1037_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block2_start_1040_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/req
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_update_start_
      -- CP-element group 293: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_sample_completed_
      -- 
    ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1040_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block2_start_1040_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1040_update_completed_
      -- 
    ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1040_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block2_start_1043_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_update_start_
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/req
      -- 
    ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1043_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block2_start_1043_inst_req_1); -- 
    -- CP-element group 296:  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (6) 
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/req
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1043_Update/$exit
      -- 
    ack_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1043_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    req_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(296), ack => WPIPE_Block2_start_1046_inst_req_0); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/req
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_update_start_
      -- CP-element group 297: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_sample_completed_
      -- 
    ack_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1046_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1046_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1046_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/$entry
      -- 
    ack_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1046_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1049_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/req
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_update_start_
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Sample/$exit
      -- 
    ack_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1049_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1049_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1049_update_completed_
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1049_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1052_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/req
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_update_start_
      -- 
    ack_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1052_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1052_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1052_Update/ack
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1052_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1055_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/req
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_update_start_
      -- CP-element group 303: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_sample_completed_
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1055_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1055_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1055_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_sample_start_
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1055_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1058_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/req
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_update_start_
      -- CP-element group 305: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_sample_completed_
      -- 
    ack_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1058_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1058_inst_req_1); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	339 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1058_update_completed_
      -- 
    ack_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1058_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	418 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/req
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_update_start_
      -- CP-element group 307: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_sample_completed_
      -- 
    ack_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1061_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block3_start_1061_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/$entry
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1061_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block3_start_1064_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_update_start_
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/req
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Sample/$exit
      -- 
    ack_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1064_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block3_start_1064_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1064_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_sample_start_
      -- 
    ack_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1064_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block3_start_1067_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/req
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_update_start_
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Sample/ack
      -- 
    ack_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1067_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block3_start_1067_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1067_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/req
      -- 
    ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1067_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block3_start_1070_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_update_start_
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/req
      -- 
    ack_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1070_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block3_start_1070_inst_req_1); -- 
    -- CP-element group 314:  transition  input  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1070_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/req
      -- 
    ack_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1070_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    req_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(314), ack => WPIPE_Block3_start_1073_inst_req_0); -- 
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_update_start_
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Sample/ack
      -- CP-element group 315: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/req
      -- 
    ack_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1073_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    req_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(315), ack => WPIPE_Block3_start_1073_inst_req_1); -- 
    -- CP-element group 316:  transition  input  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (6) 
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1073_Update/ack
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_sample_start_
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/req
      -- 
    ack_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1073_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    req_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(316), ack => WPIPE_Block3_start_1076_inst_req_0); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_update_start_
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Sample/ack
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/req
      -- 
    ack_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1076_inst_ack_0, ack => convTranspose_CP_39_elements(317)); -- 
    req_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block3_start_1076_inst_req_1); -- 
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1076_Update/ack
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/req
      -- 
    ack_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1076_inst_ack_1, ack => convTranspose_CP_39_elements(318)); -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block3_start_1079_inst_req_0); -- 
    -- CP-element group 319:  transition  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (6) 
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_update_start_
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Sample/ack
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/req
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1079_inst_ack_0, ack => convTranspose_CP_39_elements(319)); -- 
    req_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(319), ack => WPIPE_Block3_start_1079_inst_req_1); -- 
    -- CP-element group 320:  transition  input  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (6) 
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1079_Update/ack
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/req
      -- 
    ack_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1079_inst_ack_1, ack => convTranspose_CP_39_elements(320)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(320), ack => WPIPE_Block3_start_1082_inst_req_0); -- 
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_update_start_
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/req
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1082_inst_ack_0, ack => convTranspose_CP_39_elements(321)); -- 
    req_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(321), ack => WPIPE_Block3_start_1082_inst_req_1); -- 
    -- CP-element group 322:  transition  input  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (6) 
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1082_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/req
      -- 
    ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1082_inst_ack_1, ack => convTranspose_CP_39_elements(322)); -- 
    req_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block3_start_1085_inst_req_0); -- 
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_update_start_
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/req
      -- 
    ack_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1085_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block3_start_1085_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1085_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/req
      -- 
    ack_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1085_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block3_start_1088_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_update_start_
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/req
      -- 
    ack_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1088_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block3_start_1088_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1088_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/req
      -- 
    ack_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1088_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block3_start_1091_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_update_start_
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/req
      -- 
    ack_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1091_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block3_start_1091_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1091_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/req
      -- 
    ack_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1091_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block3_start_1094_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_update_start_
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/req
      -- 
    ack_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1094_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block3_start_1094_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	339 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1094_Update/ack
      -- 
    ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1094_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	418 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_update_start_
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/ra
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/cr
      -- 
    ra_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1098_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    cr_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => RPIPE_Block0_done_1098_inst_req_1); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	339 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Update/ca
      -- 
    ca_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1098_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	418 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_update_start_
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/ra
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/cr
      -- 
    ra_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1101_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    cr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => RPIPE_Block1_done_1101_inst_req_1); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	339 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Update/ca
      -- 
    ca_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1101_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	418 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_update_start_
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/ra
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/cr
      -- 
    ra_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1104_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    cr_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => RPIPE_Block2_done_1104_inst_req_1); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	339 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Update/ca
      -- 
    ca_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1104_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	418 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_update_start_
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/ra
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/cr
      -- 
    ra_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1107_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    cr_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => RPIPE_Block3_done_1107_inst_req_1); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Update/ca
      -- 
    ca_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1107_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    -- CP-element group 339:  join  fork  transition  place  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	282 
    -- CP-element group 339: 	306 
    -- CP-element group 339: 	330 
    -- CP-element group 339: 	332 
    -- CP-element group 339: 	334 
    -- CP-element group 339: 	336 
    -- CP-element group 339: 	338 
    -- CP-element group 339: 	234 
    -- CP-element group 339: 	258 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339: 	341 
    -- CP-element group 339: 	343 
    -- CP-element group 339:  members (13) 
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108__exit__
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124__entry__
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/$exit
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_update_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/crr
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/ccr
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_update_start_
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/cr
      -- 
    crr_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => call_stmt_1111_call_req_0); -- 
    ccr_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => call_stmt_1111_call_req_1); -- 
    cr_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => type_cast_1115_inst_req_1); -- 
    convTranspose_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(282) & convTranspose_CP_39_elements(306) & convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(332) & convTranspose_CP_39_elements(334) & convTranspose_CP_39_elements(336) & convTranspose_CP_39_elements(338) & convTranspose_CP_39_elements(234) & convTranspose_CP_39_elements(258);
      gj_convTranspose_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Sample/cra
      -- 
    cra_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1111_call_ack_0, ack => convTranspose_CP_39_elements(340)); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/call_stmt_1111_Update/cca
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/rr
      -- 
    cca_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1111_call_ack_1, ack => convTranspose_CP_39_elements(341)); -- 
    rr_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => type_cast_1115_inst_req_0); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_sample_completed_
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Sample/ra
      -- 
    ra_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_0, ack => convTranspose_CP_39_elements(342)); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	339 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_update_completed_
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/type_cast_1115_Update/ca
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_sample_start_
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/req
      -- 
    ca_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1115_inst_ack_1, ack => convTranspose_CP_39_elements(343)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_elapsed_time_pipe_1122_inst_req_0); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_sample_completed_
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_update_start_
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Sample/ack
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/req
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1122_inst_ack_0, ack => convTranspose_CP_39_elements(344)); -- 
    req_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_elapsed_time_pipe_1122_inst_req_1); -- 
    -- CP-element group 345:  branch  transition  place  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (17) 
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124__exit__
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_1131__entry__
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_1131__exit__
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132__entry__
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_update_completed_
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/call_stmt_1111_to_assign_stmt_1124/WPIPE_elapsed_time_pipe_1122_Update/ack
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_1131/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/assign_stmt_1131/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132_dead_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132_eval_test/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132_eval_test/$exit
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132_eval_test/branch_req
      -- CP-element group 345: 	 branch_block_stmt_33/R_cmp330406_1133_place
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132_if_link/$entry
      -- CP-element group 345: 	 branch_block_stmt_33/if_stmt_1132_else_link/$entry
      -- 
    ack_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1122_inst_ack_1, ack => convTranspose_CP_39_elements(345)); -- 
    branch_req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => if_stmt_1132_branch_req_0); -- 
    -- CP-element group 346:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: 	349 
    -- CP-element group 346:  members (18) 
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1138__exit__
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173__entry__
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1138_PhiReqMerge
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1138_PhiAck/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1138_PhiAck/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend259_bbx_xnph_PhiReq/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/if_stmt_1132_if_link/$exit
      -- CP-element group 346: 	 branch_block_stmt_33/if_stmt_1132_if_link/if_choice_transition
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend259_bbx_xnph
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_33/forx_xend259_bbx_xnph_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_update_start_
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Sample/rr
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Update/cr
      -- CP-element group 346: 	 branch_block_stmt_33/merge_stmt_1138_PhiAck/dummy
      -- 
    if_choice_transition_2675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1132_branch_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    rr_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => type_cast_1159_inst_req_0); -- 
    cr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => type_cast_1159_inst_req_1); -- 
    -- CP-element group 347:  transition  place  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	425 
    -- CP-element group 347:  members (5) 
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xend259_forx_xend404_PhiReq/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xend259_forx_xend404_PhiReq/$entry
      -- CP-element group 347: 	 branch_block_stmt_33/if_stmt_1132_else_link/$exit
      -- CP-element group 347: 	 branch_block_stmt_33/if_stmt_1132_else_link/else_choice_transition
      -- CP-element group 347: 	 branch_block_stmt_33/forx_xend259_forx_xend404
      -- 
    else_choice_transition_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1132_branch_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Sample/ra
      -- 
    ra_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_0, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  place  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	346 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	419 
    -- CP-element group 349:  members (9) 
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173__exit__
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_33/assign_stmt_1144_to_assign_stmt_1173/type_cast_1159_Update/ca
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/$entry
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1176/$entry
      -- CP-element group 349: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/$entry
      -- 
    ca_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_1, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	424 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	395 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_sample_complete
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Sample/ack
      -- 
    ack_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1188_index_offset_ack_0, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  transition  input  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	424 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (11) 
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_root_address_calculated
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_offset_calculated
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Update/ack
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_base_plus_offset/$entry
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_base_plus_offset/$exit
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_base_plus_offset/sum_rename_req
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_base_plus_offset/sum_rename_ack
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_request/$entry
      -- CP-element group 351: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_request/req
      -- 
    ack_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1188_index_offset_ack_1, ack => convTranspose_CP_39_elements(351)); -- 
    req_2741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => addr_of_1189_final_reg_req_0); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_request/$exit
      -- CP-element group 352: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_request/ack
      -- 
    ack_2742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1189_final_reg_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    -- CP-element group 353:  join  fork  transition  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	424 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (24) 
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_complete/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_complete/ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_word_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_address_resized
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_addr_resize/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_addr_resize/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_addr_resize/base_resize_req
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_addr_resize/base_resize_ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_plus_offset/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_plus_offset/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_plus_offset/sum_rename_req
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_base_plus_offset/sum_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_word_addrgen/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_word_addrgen/$exit
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_word_addrgen/root_register_req
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_word_addrgen/root_register_ack
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/word_access_start/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/word_access_start/word_0/$entry
      -- CP-element group 353: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/word_access_start/word_0/rr
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1189_final_reg_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    rr_2780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(353), ack => ptr_deref_1193_load_0_req_0); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (5) 
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/word_access_start/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/word_access_start/word_0/$exit
      -- CP-element group 354: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Sample/word_access_start/word_0/ra
      -- 
    ra_2781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1193_load_0_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  fork  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	424 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355: 	358 
    -- CP-element group 355: 	360 
    -- CP-element group 355: 	362 
    -- CP-element group 355: 	364 
    -- CP-element group 355: 	366 
    -- CP-element group 355: 	368 
    -- CP-element group 355: 	370 
    -- CP-element group 355:  members (33) 
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/word_access_complete/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/word_access_complete/word_0/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/word_access_complete/word_0/ca
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/ptr_deref_1193_Merge/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/ptr_deref_1193_Merge/$exit
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/ptr_deref_1193_Merge/merge_req
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/ptr_deref_1193_Merge/merge_ack
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_sample_start_
      -- 
    ca_2792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1193_load_0_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    rr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1197_inst_req_0); -- 
    rr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1207_inst_req_0); -- 
    rr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1217_inst_req_0); -- 
    rr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1227_inst_req_0); -- 
    rr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1237_inst_req_0); -- 
    rr_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1247_inst_req_0); -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1257_inst_req_0); -- 
    rr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => type_cast_1267_inst_req_0); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Sample/ra
      -- 
    ra_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_0, ack => convTranspose_CP_39_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	424 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	392 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Update/ca
      -- 
    ca_2811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_1, ack => convTranspose_CP_39_elements(357)); -- 
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	355 
    -- CP-element group 358: successors 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_sample_completed_
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Sample/ra
      -- 
    ra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_0, ack => convTranspose_CP_39_elements(358)); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	424 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	389 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Update/ca
      -- 
    ca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_1, ack => convTranspose_CP_39_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	355 
    -- CP-element group 360: successors 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Sample/ra
      -- 
    ra_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1217_inst_ack_0, ack => convTranspose_CP_39_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	424 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	386 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Update/ca
      -- 
    ca_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1217_inst_ack_1, ack => convTranspose_CP_39_elements(361)); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	355 
    -- CP-element group 362: successors 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Sample/ra
      -- 
    ra_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_0, ack => convTranspose_CP_39_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	424 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	383 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Update/ca
      -- 
    ca_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_1, ack => convTranspose_CP_39_elements(363)); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	355 
    -- CP-element group 364: successors 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Sample/ra
      -- 
    ra_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1237_inst_ack_0, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	424 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	380 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Update/ca
      -- 
    ca_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1237_inst_ack_1, ack => convTranspose_CP_39_elements(365)); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	355 
    -- CP-element group 366: successors 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Sample/ra
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_sample_completed_
      -- 
    ra_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_0, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	424 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	377 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Update/ca
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_update_completed_
      -- 
    ca_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1247_inst_ack_1, ack => convTranspose_CP_39_elements(367)); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	355 
    -- CP-element group 368: successors 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Sample/ra
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1257_inst_ack_0, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	424 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Update/ca
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1257_inst_ack_1, ack => convTranspose_CP_39_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	355 
    -- CP-element group 370: successors 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Sample/ra
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_sample_completed_
      -- 
    ra_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1267_inst_ack_0, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	424 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Update/ca
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Sample/req
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_update_completed_
      -- 
    ca_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1267_inst_ack_1, ack => convTranspose_CP_39_elements(371)); -- 
    req_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => WPIPE_ConvTranspose_output_pipe_1269_inst_req_0); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Update/req
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Sample/ack
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_update_start_
      -- CP-element group 372: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_sample_completed_
      -- 
    ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1269_inst_ack_0, ack => convTranspose_CP_39_elements(372)); -- 
    req_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => WPIPE_ConvTranspose_output_pipe_1269_inst_req_1); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Update/ack
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1269_update_completed_
      -- 
    ack_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1269_inst_ack_1, ack => convTranspose_CP_39_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Sample/req
      -- CP-element group 374: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_sample_start_
      -- 
    req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(374), ack => WPIPE_ConvTranspose_output_pipe_1272_inst_req_0); -- 
    convTranspose_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(369) & convTranspose_CP_39_elements(373);
      gj_convTranspose_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Sample/ack
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Update/req
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_update_start_
      -- CP-element group 375: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_sample_completed_
      -- 
    ack_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1272_inst_ack_0, ack => convTranspose_CP_39_elements(375)); -- 
    req_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => WPIPE_ConvTranspose_output_pipe_1272_inst_req_1); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_Update/ack
      -- CP-element group 376: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1272_update_completed_
      -- 
    ack_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1272_inst_ack_1, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	367 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Sample/req
      -- CP-element group 377: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Sample/$entry
      -- 
    req_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => WPIPE_ConvTranspose_output_pipe_1275_inst_req_0); -- 
    convTranspose_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(367) & convTranspose_CP_39_elements(376);
      gj_convTranspose_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Update/req
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_update_start_
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Sample/$exit
      -- 
    ack_2946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1275_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    req_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => WPIPE_ConvTranspose_output_pipe_1275_inst_req_1); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1275_Update/ack
      -- 
    ack_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1275_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	365 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Sample/req
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_sample_start_
      -- 
    req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => WPIPE_ConvTranspose_output_pipe_1278_inst_req_0); -- 
    convTranspose_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(365) & convTranspose_CP_39_elements(379);
      gj_convTranspose_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (6) 
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Update/req
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Update/$entry
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Sample/ack
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_update_start_
      -- CP-element group 381: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_sample_completed_
      -- 
    ack_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1278_inst_ack_0, ack => convTranspose_CP_39_elements(381)); -- 
    req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(381), ack => WPIPE_ConvTranspose_output_pipe_1278_inst_req_1); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Update/ack
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1278_update_completed_
      -- 
    ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1278_inst_ack_1, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	363 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Sample/req
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_sample_start_
      -- 
    req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(383), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_0); -- 
    convTranspose_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(363) & convTranspose_CP_39_elements(382);
      gj_convTranspose_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  transition  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Update/req
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Sample/ack
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_update_start_
      -- CP-element group 384: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_sample_completed_
      -- 
    ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => WPIPE_ConvTranspose_output_pipe_1281_inst_req_1); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Update/ack
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1281_update_completed_
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    -- CP-element group 386:  join  transition  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	361 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Sample/req
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Sample/$entry
      -- CP-element group 386: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_sample_start_
      -- 
    req_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_0); -- 
    convTranspose_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(361) & convTranspose_CP_39_elements(385);
      gj_convTranspose_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (6) 
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Update/req
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Sample/ack
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_update_start_
      -- CP-element group 387: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_sample_completed_
      -- 
    ack_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0, ack => convTranspose_CP_39_elements(387)); -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(387), ack => WPIPE_ConvTranspose_output_pipe_1284_inst_req_1); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Update/ack
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1284_update_completed_
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1, ack => convTranspose_CP_39_elements(388)); -- 
    -- CP-element group 389:  join  transition  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	359 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Sample/req
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Sample/$entry
      -- 
    req_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_0); -- 
    convTranspose_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(359) & convTranspose_CP_39_elements(388);
      gj_convTranspose_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_update_start_
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Update/req
      -- 
    ack_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_1); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1287_Update/ack
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    -- CP-element group 392:  join  transition  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	357 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_sample_start_
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Sample/$entry
      -- CP-element group 392: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Sample/req
      -- 
    req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(392), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_0); -- 
    convTranspose_cp_element_group_392: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_392"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(357) & convTranspose_CP_39_elements(391);
      gj_convTranspose_cp_element_group_392 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(392), clk => clk, reset => reset); --
    end block;
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_update_start_
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Update/req
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Sample/ack
      -- CP-element group 393: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Sample/$exit
      -- 
    ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0, ack => convTranspose_CP_39_elements(393)); -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(393), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_1); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Update/ack
      -- CP-element group 394: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1290_Update/$exit
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1, ack => convTranspose_CP_39_elements(394)); -- 
    -- CP-element group 395:  branch  join  transition  place  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	350 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (10) 
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303__exit__
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304__entry__
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304_else_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304_if_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304_eval_test/branch_req
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304_eval_test/$exit
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304_eval_test/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/R_exitcond1_1305_place
      -- CP-element group 395: 	 branch_block_stmt_33/if_stmt_1304_dead_link/$entry
      -- CP-element group 395: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/$exit
      -- 
    branch_req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => if_stmt_1304_branch_req_0); -- 
    convTranspose_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(350) & convTranspose_CP_39_elements(394);
      gj_convTranspose_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  merge  transition  place  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	425 
    -- CP-element group 396:  members (13) 
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1310__exit__
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xend404x_xloopexit_forx_xend404
      -- CP-element group 396: 	 branch_block_stmt_33/if_stmt_1304_if_link/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/if_stmt_1304_if_link/if_choice_transition
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1310_PhiAck/dummy
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1310_PhiAck/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1310_PhiAck/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/merge_stmt_1310_PhiReqMerge
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xbody332_forx_xend404x_xloopexit_PhiReq/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xbody332_forx_xend404x_xloopexit_PhiReq/$entry
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xbody332_forx_xend404x_xloopexit
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xend404x_xloopexit_forx_xend404_PhiReq/$exit
      -- CP-element group 396: 	 branch_block_stmt_33/forx_xend404x_xloopexit_forx_xend404_PhiReq/$entry
      -- 
    if_choice_transition_3034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1304_branch_ack_1, ack => convTranspose_CP_39_elements(396)); -- 
    -- CP-element group 397:  fork  transition  place  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	420 
    -- CP-element group 397: 	421 
    -- CP-element group 397:  members (12) 
      -- CP-element group 397: 	 branch_block_stmt_33/if_stmt_1304_else_link/$exit
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/if_stmt_1304_else_link/else_choice_transition
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Update/cr
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Sample/rr
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/$entry
      -- CP-element group 397: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/$entry
      -- 
    else_choice_transition_3038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1304_branch_ack_0, ack => convTranspose_CP_39_elements(397)); -- 
    cr_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => type_cast_1179_inst_req_1); -- 
    rr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => type_cast_1179_inst_req_0); -- 
    -- CP-element group 398:  merge  branch  transition  place  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	165 
    -- CP-element group 398: 	120 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	121 
    -- CP-element group 398: 	122 
    -- CP-element group 398:  members (17) 
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402__exit__
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408__entry__
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408__exit__
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409__entry__
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/assign_stmt_408/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_dead_link/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_eval_test/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_eval_test/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_eval_test/branch_req
      -- CP-element group 398: 	 branch_block_stmt_33/R_cmp180413_410_place
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_if_link/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/if_stmt_409_else_link/$entry
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiReqMerge
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiAck/dummy
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiAck/$exit
      -- CP-element group 398: 	 branch_block_stmt_33/merge_stmt_402_PhiAck/$entry
      -- 
    branch_req_927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => if_stmt_409_branch_req_0); -- 
    convTranspose_CP_39_elements(398) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 399:  transition  output  delay-element  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	124 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	403 
    -- CP-element group 399:  members (5) 
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_req
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_457_konst_delay_trans
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$exit
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/phi_stmt_453/$exit
      -- CP-element group 399: 	 branch_block_stmt_33/bbx_xnph419_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_453_req_3086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_req_3086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => phi_stmt_453_req_0); -- 
    -- Element group convTranspose_CP_39_elements(399) is a control-delay.
    cp_element_399_delay: control_delay_element  generic map(name => " 399_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(399), clk => clk, reset =>reset);
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	166 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	402 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/ra
      -- CP-element group 400: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Sample/$exit
      -- 
    ra_3106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_459_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	166 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (2) 
      -- CP-element group 401: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/ca
      -- CP-element group 401: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/Update/$exit
      -- 
    ca_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_459_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	400 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_req
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/SplitProtocol/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/type_cast_459/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/phi_stmt_453_sources/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/phi_stmt_453/$exit
      -- CP-element group 402: 	 branch_block_stmt_33/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_453_req_3112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_req_3112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => phi_stmt_453_req_1); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(400) & convTranspose_CP_39_elements(401);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  merge  transition  place  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	399 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_33/merge_stmt_452_PhiReqMerge
      -- CP-element group 403: 	 branch_block_stmt_33/merge_stmt_452_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(403) <= OrReduce(convTranspose_CP_39_elements(399) & convTranspose_CP_39_elements(402));
    -- CP-element group 404:  fork  transition  place  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	160 
    -- CP-element group 404: 	163 
    -- CP-element group 404: 	125 
    -- CP-element group 404: 	126 
    -- CP-element group 404: 	128 
    -- CP-element group 404: 	129 
    -- CP-element group 404: 	132 
    -- CP-element group 404: 	136 
    -- CP-element group 404: 	140 
    -- CP-element group 404: 	144 
    -- CP-element group 404: 	148 
    -- CP-element group 404: 	152 
    -- CP-element group 404: 	156 
    -- CP-element group 404:  members (56) 
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/merge_stmt_452__exit__
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615__entry__
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_558_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_540_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/word_0/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/word_access_complete/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_522_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_576_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_594_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/ptr_deref_602_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resized_1
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scaled_1
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_computed_1
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/index_resize_req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_resize_1/index_resize_ack
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/$exit
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/scale_rename_req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_index_scale_1/scale_rename_ack
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_update_start
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Sample/req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/array_obj_ref_465_final_index_sum_regn_Update/req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/addr_of_466_complete/req
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_sample_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/RPIPE_ConvTranspose_input_pipe_469_Sample/rr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_473_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_486_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_33/assign_stmt_467_to_assign_stmt_615/type_cast_504_update_start_
      -- CP-element group 404: 	 branch_block_stmt_33/merge_stmt_452_PhiAck/phi_stmt_453_ack
      -- CP-element group 404: 	 branch_block_stmt_33/merge_stmt_452_PhiAck/$exit
      -- 
    phi_stmt_453_ack_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_453_ack_0, ack => convTranspose_CP_39_elements(404)); -- 
    cr_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_558_inst_req_1); -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_540_inst_req_1); -- 
    cr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_504_inst_req_1); -- 
    cr_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => ptr_deref_602_store_0_req_1); -- 
    cr_1199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_576_inst_req_1); -- 
    cr_1115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_522_inst_req_1); -- 
    cr_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_594_inst_req_1); -- 
    req_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => array_obj_ref_465_index_offset_req_0); -- 
    req_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => array_obj_ref_465_index_offset_req_1); -- 
    req_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => addr_of_466_final_reg_req_1); -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => RPIPE_ConvTranspose_input_pipe_469_inst_req_0); -- 
    cr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_473_inst_req_1); -- 
    cr_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_486_inst_req_1); -- 
    -- CP-element group 405:  transition  output  delay-element  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	168 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	409 
    -- CP-element group 405:  members (5) 
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_666_konst_delay_trans
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$exit
      -- CP-element group 405: 	 branch_block_stmt_33/bbx_xnph415_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_req
      -- 
    phi_stmt_660_req_3140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_660_req_3140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => phi_stmt_660_req_1); -- 
    -- Element group convTranspose_CP_39_elements(405) is a control-delay.
    cp_element_405_delay: control_delay_element  generic map(name => " 405_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(405), clk => clk, reset =>reset);
    -- CP-element group 406:  transition  input  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	210 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/ra
      -- CP-element group 406: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Sample/$exit
      -- 
    ra_3160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_663_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	210 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (2) 
      -- CP-element group 407: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/ca
      -- CP-element group 407: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/Update/$exit
      -- 
    ca_3165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_663_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (6) 
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_req
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/SplitProtocol/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/type_cast_663/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/phi_stmt_660_sources/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/phi_stmt_660/$exit
      -- CP-element group 408: 	 branch_block_stmt_33/forx_xbody182_forx_xbody182_PhiReq/$exit
      -- 
    phi_stmt_660_req_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_660_req_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => phi_stmt_660_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(406) & convTranspose_CP_39_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  merge  transition  place  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	405 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (2) 
      -- CP-element group 409: 	 branch_block_stmt_33/merge_stmt_659_PhiReqMerge
      -- CP-element group 409: 	 branch_block_stmt_33/merge_stmt_659_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(409) <= OrReduce(convTranspose_CP_39_elements(405) & convTranspose_CP_39_elements(408));
    -- CP-element group 410:  fork  transition  place  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	180 
    -- CP-element group 410: 	184 
    -- CP-element group 410: 	188 
    -- CP-element group 410: 	192 
    -- CP-element group 410: 	196 
    -- CP-element group 410: 	200 
    -- CP-element group 410: 	204 
    -- CP-element group 410: 	207 
    -- CP-element group 410: 	172 
    -- CP-element group 410: 	173 
    -- CP-element group 410: 	176 
    -- CP-element group 410: 	169 
    -- CP-element group 410: 	170 
    -- CP-element group 410:  members (56) 
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_sample_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/merge_stmt_659__exit__
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822__entry__
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/scale_rename_ack
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/scale_rename_req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/$exit
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scale_1/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/index_resize_ack
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/index_resize_req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_complete/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/req
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/$exit
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_680_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resize_1/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_computed_1
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_scaled_1
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_index_resized_1
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_711_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/array_obj_ref_672_final_index_sum_regn_update_start
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/addr_of_673_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/rr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/RPIPE_ConvTranspose_input_pipe_676_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_693_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_729_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_747_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_765_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_783_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/type_cast_801_Update/cr
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_update_start_
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/$entry
      -- CP-element group 410: 	 branch_block_stmt_33/assign_stmt_674_to_assign_stmt_822/ptr_deref_809_Update/word_access_complete/word_0/cr
      -- CP-element group 410: 	 branch_block_stmt_33/merge_stmt_659_PhiAck/phi_stmt_660_ack
      -- CP-element group 410: 	 branch_block_stmt_33/merge_stmt_659_PhiAck/$exit
      -- 
    phi_stmt_660_ack_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_660_ack_0, ack => convTranspose_CP_39_elements(410)); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_711_inst_req_1); -- 
    req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => array_obj_ref_672_index_offset_req_1); -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_693_inst_req_1); -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_680_inst_req_1); -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => addr_of_673_final_reg_req_1); -- 
    req_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => array_obj_ref_672_index_offset_req_0); -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => RPIPE_ConvTranspose_input_pipe_676_inst_req_0); -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_729_inst_req_1); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_747_inst_req_1); -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_765_inst_req_1); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_783_inst_req_1); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => type_cast_801_inst_req_1); -- 
    cr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => ptr_deref_809_store_0_req_1); -- 
    -- CP-element group 411:  merge  fork  transition  place  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	209 
    -- CP-element group 411: 	122 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	211 
    -- CP-element group 411: 	212 
    -- CP-element group 411: 	213 
    -- CP-element group 411: 	214 
    -- CP-element group 411: 	215 
    -- CP-element group 411: 	216 
    -- CP-element group 411:  members (25) 
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831__exit__
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859__entry__
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiReqMerge
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Sample/rr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_834_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Sample/rr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_838_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_update_start_
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Sample/rr
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_33/assign_stmt_835_to_assign_stmt_859/type_cast_842_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiAck/dummy
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiAck/$exit
      -- CP-element group 411: 	 branch_block_stmt_33/merge_stmt_831_PhiAck/$entry
      -- 
    rr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_834_inst_req_0); -- 
    cr_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_834_inst_req_1); -- 
    rr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_838_inst_req_0); -- 
    cr_1686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_838_inst_req_1); -- 
    rr_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_842_inst_req_0); -- 
    cr_1700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => type_cast_842_inst_req_1); -- 
    convTranspose_CP_39_elements(411) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 412:  transition  output  delay-element  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	221 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	416 
    -- CP-element group 412:  members (5) 
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$exit
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_908_konst_delay_trans
      -- CP-element group 412: 	 branch_block_stmt_33/bbx_xnph411_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_req
      -- 
    phi_stmt_904_req_3217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_904_req_3217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => phi_stmt_904_req_0); -- 
    -- Element group convTranspose_CP_39_elements(412) is a control-delay.
    cp_element_412_delay: control_delay_element  generic map(name => " 412_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(412), clk => clk, reset =>reset);
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	230 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	415 
    -- CP-element group 413:  members (2) 
      -- CP-element group 413: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/ra
      -- CP-element group 413: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Sample/$exit
      -- 
    ra_3237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_910_inst_ack_0, ack => convTranspose_CP_39_elements(413)); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	230 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (2) 
      -- CP-element group 414: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/ca
      -- CP-element group 414: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/Update/$exit
      -- 
    ca_3242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_910_inst_ack_1, ack => convTranspose_CP_39_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	413 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_req
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/SplitProtocol/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/type_cast_910/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/phi_stmt_904_sources/$exit
      -- CP-element group 415: 	 branch_block_stmt_33/forx_xbody252_forx_xbody252_PhiReq/phi_stmt_904/$exit
      -- 
    phi_stmt_904_req_3243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_904_req_3243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => phi_stmt_904_req_1); -- 
    convTranspose_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(413) & convTranspose_CP_39_elements(414);
      gj_convTranspose_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  merge  transition  place  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	412 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (2) 
      -- CP-element group 416: 	 branch_block_stmt_33/merge_stmt_903_PhiReqMerge
      -- CP-element group 416: 	 branch_block_stmt_33/merge_stmt_903_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(416) <= OrReduce(convTranspose_CP_39_elements(412) & convTranspose_CP_39_elements(415));
    -- CP-element group 417:  fork  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	222 
    -- CP-element group 417: 	223 
    -- CP-element group 417: 	225 
    -- CP-element group 417: 	227 
    -- CP-element group 417:  members (29) 
      -- CP-element group 417: 	 branch_block_stmt_33/merge_stmt_903_PhiAck/phi_stmt_904_ack
      -- CP-element group 417: 	 branch_block_stmt_33/merge_stmt_903__exit__
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934__entry__
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_update_start_
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resized_1
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scaled_1
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_computed_1
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/$exit
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/index_resize_req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_resize_1/index_resize_ack
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/$exit
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/scale_rename_req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_index_scale_1/scale_rename_ack
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_update_start
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Sample/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/array_obj_ref_916_final_index_sum_regn_Update/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/addr_of_917_complete/req
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_update_start_
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/$entry
      -- CP-element group 417: 	 branch_block_stmt_33/assign_stmt_918_to_assign_stmt_934/ptr_deref_920_Update/word_access_complete/word_0/cr
      -- CP-element group 417: 	 branch_block_stmt_33/merge_stmt_903_PhiAck/$exit
      -- 
    phi_stmt_904_ack_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_904_ack_0, ack => convTranspose_CP_39_elements(417)); -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => array_obj_ref_916_index_offset_req_0); -- 
    req_1770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => array_obj_ref_916_index_offset_req_1); -- 
    req_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => addr_of_917_final_reg_req_1); -- 
    cr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => ptr_deref_920_store_0_req_1); -- 
    -- CP-element group 418:  merge  fork  transition  place  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	219 
    -- CP-element group 418: 	229 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	283 
    -- CP-element group 418: 	307 
    -- CP-element group 418: 	331 
    -- CP-element group 418: 	333 
    -- CP-element group 418: 	335 
    -- CP-element group 418: 	337 
    -- CP-element group 418: 	231 
    -- CP-element group 418: 	232 
    -- CP-element group 418: 	234 
    -- CP-element group 418: 	235 
    -- CP-element group 418: 	259 
    -- CP-element group 418:  members (40) 
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943__exit__
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108__entry__
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiReqMerge
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block3_start_1061_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/$exit
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block1_start_989_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block2_start_1025_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_update_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Sample/crr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/call_stmt_946_Update/ccr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_update_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/type_cast_951_Update/cr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/WPIPE_Block0_start_953_Sample/req
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block0_done_1098_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block1_done_1101_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block2_done_1104_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_33/call_stmt_946_to_assign_stmt_1108/RPIPE_Block3_done_1107_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_33/merge_stmt_943_PhiAck/dummy
      -- 
    req_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block3_start_1061_inst_req_0); -- 
    req_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block1_start_989_inst_req_0); -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block2_start_1025_inst_req_0); -- 
    crr_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => call_stmt_946_call_req_0); -- 
    ccr_1871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => call_stmt_946_call_req_1); -- 
    cr_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => type_cast_951_inst_req_1); -- 
    req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => WPIPE_Block0_start_953_inst_req_0); -- 
    rr_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block0_done_1098_inst_req_0); -- 
    rr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block1_done_1101_inst_req_0); -- 
    rr_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block2_done_1104_inst_req_0); -- 
    rr_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(418), ack => RPIPE_Block3_done_1107_inst_req_0); -- 
    convTranspose_CP_39_elements(418) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 419:  transition  output  delay-element  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	349 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	423 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_req
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1182_konst_delay_trans
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/phi_stmt_1176/$exit
      -- CP-element group 419: 	 branch_block_stmt_33/bbx_xnph_forx_xbody332_PhiReq/$exit
      -- 
    phi_stmt_1176_req_3294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1176_req_3294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(419), ack => phi_stmt_1176_req_1); -- 
    -- Element group convTranspose_CP_39_elements(419) is a control-delay.
    cp_element_419_delay: control_delay_element  generic map(name => " 419_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(349), ack => convTranspose_CP_39_elements(419), clk => clk, reset =>reset);
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	397 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	422 
    -- CP-element group 420:  members (2) 
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Sample/ra
      -- CP-element group 420: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Sample/$exit
      -- 
    ra_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_0, ack => convTranspose_CP_39_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	397 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (2) 
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Update/ca
      -- CP-element group 421: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/Update/$exit
      -- 
    ca_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_1, ack => convTranspose_CP_39_elements(421)); -- 
    -- CP-element group 422:  join  transition  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (6) 
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/SplitProtocol/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/type_cast_1179/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_req
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/phi_stmt_1176_sources/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/phi_stmt_1176/$exit
      -- CP-element group 422: 	 branch_block_stmt_33/forx_xbody332_forx_xbody332_PhiReq/$exit
      -- 
    phi_stmt_1176_req_3320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1176_req_3320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(422), ack => phi_stmt_1176_req_0); -- 
    convTranspose_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(420) & convTranspose_CP_39_elements(421);
      gj_convTranspose_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  merge  transition  place  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	419 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (2) 
      -- CP-element group 423: 	 branch_block_stmt_33/merge_stmt_1175_PhiAck/$entry
      -- CP-element group 423: 	 branch_block_stmt_33/merge_stmt_1175_PhiReqMerge
      -- 
    convTranspose_CP_39_elements(423) <= OrReduce(convTranspose_CP_39_elements(419) & convTranspose_CP_39_elements(422));
    -- CP-element group 424:  fork  transition  place  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	350 
    -- CP-element group 424: 	351 
    -- CP-element group 424: 	353 
    -- CP-element group 424: 	355 
    -- CP-element group 424: 	357 
    -- CP-element group 424: 	359 
    -- CP-element group 424: 	361 
    -- CP-element group 424: 	363 
    -- CP-element group 424: 	365 
    -- CP-element group 424: 	367 
    -- CP-element group 424: 	369 
    -- CP-element group 424: 	371 
    -- CP-element group 424:  members (53) 
      -- CP-element group 424: 	 branch_block_stmt_33/merge_stmt_1175__exit__
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303__entry__
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/merge_stmt_1175_PhiAck/phi_stmt_1176_ack
      -- CP-element group 424: 	 branch_block_stmt_33/merge_stmt_1175_PhiAck/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1267_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_resized_1
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_scaled_1
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_computed_1
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_resize_1/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_resize_1/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_resize_1/index_resize_req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_resize_1/index_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_scale_1/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_scale_1/$exit
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_scale_1/scale_rename_req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_index_scale_1/scale_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_update_start
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Sample/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/array_obj_ref_1188_final_index_sum_regn_Update/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/addr_of_1189_complete/req
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1257_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/word_access_complete/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/word_access_complete/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/ptr_deref_1193_Update/word_access_complete/word_0/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1197_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1207_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1217_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1227_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_update_start_
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1237_Update/cr
      -- CP-element group 424: 	 branch_block_stmt_33/assign_stmt_1190_to_assign_stmt_1303/type_cast_1247_update_start_
      -- 
    phi_stmt_1176_ack_3325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1176_ack_0, ack => convTranspose_CP_39_elements(424)); -- 
    cr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1267_inst_req_1); -- 
    cr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1247_inst_req_1); -- 
    req_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => array_obj_ref_1188_index_offset_req_0); -- 
    req_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => array_obj_ref_1188_index_offset_req_1); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => addr_of_1189_final_reg_req_1); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1257_inst_req_1); -- 
    cr_2791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => ptr_deref_1193_load_0_req_1); -- 
    cr_2810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1197_inst_req_1); -- 
    cr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1207_inst_req_1); -- 
    cr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1217_inst_req_1); -- 
    cr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1227_inst_req_1); -- 
    cr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => type_cast_1237_inst_req_1); -- 
    -- CP-element group 425:  merge  transition  place  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	347 
    -- CP-element group 425: 	396 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (16) 
      -- CP-element group 425: 	 $exit
      -- CP-element group 425: 	 branch_block_stmt_33/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/branch_block_stmt_33__exit__
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1312__exit__
      -- CP-element group 425: 	 branch_block_stmt_33/return__
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1314__exit__
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1314_PhiAck/dummy
      -- CP-element group 425: 	 branch_block_stmt_33/return___PhiReq/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/return___PhiReq/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1314_PhiAck/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1314_PhiAck/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1314_PhiReqMerge
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1312_PhiAck/dummy
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1312_PhiAck/$exit
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1312_PhiAck/$entry
      -- CP-element group 425: 	 branch_block_stmt_33/merge_stmt_1312_PhiReqMerge
      -- 
    convTranspose_CP_39_elements(425) <= OrReduce(convTranspose_CP_39_elements(347) & convTranspose_CP_39_elements(396));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar429_915_resized : std_logic_vector(13 downto 0);
    signal R_indvar429_915_scaled : std_logic_vector(13 downto 0);
    signal R_indvar443_671_resized : std_logic_vector(10 downto 0);
    signal R_indvar443_671_scaled : std_logic_vector(10 downto 0);
    signal R_indvar459_464_resized : std_logic_vector(13 downto 0);
    signal R_indvar459_464_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1187_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1187_scaled : std_logic_vector(13 downto 0);
    signal add104_336 : std_logic_vector(15 downto 0);
    signal add113_361 : std_logic_vector(15 downto 0);
    signal add122_386 : std_logic_vector(15 downto 0);
    signal add12_83 : std_logic_vector(15 downto 0);
    signal add136_492 : std_logic_vector(63 downto 0);
    signal add142_510 : std_logic_vector(63 downto 0);
    signal add148_528 : std_logic_vector(63 downto 0);
    signal add154_546 : std_logic_vector(63 downto 0);
    signal add160_564 : std_logic_vector(63 downto 0);
    signal add166_582 : std_logic_vector(63 downto 0);
    signal add172_600 : std_logic_vector(63 downto 0);
    signal add192_699 : std_logic_vector(63 downto 0);
    signal add198_717 : std_logic_vector(63 downto 0);
    signal add204_735 : std_logic_vector(63 downto 0);
    signal add210_753 : std_logic_vector(63 downto 0);
    signal add216_771 : std_logic_vector(63 downto 0);
    signal add21_108 : std_logic_vector(15 downto 0);
    signal add222_789 : std_logic_vector(63 downto 0);
    signal add228_807 : std_logic_vector(63 downto 0);
    signal add30_133 : std_logic_vector(15 downto 0);
    signal add39_158 : std_logic_vector(15 downto 0);
    signal add48_183 : std_logic_vector(15 downto 0);
    signal add57_208 : std_logic_vector(15 downto 0);
    signal add86_286 : std_logic_vector(15 downto 0);
    signal add95_311 : std_logic_vector(15 downto 0);
    signal add_58 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1188_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1188_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1188_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1188_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1188_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1188_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_465_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_672_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_672_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_916_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_916_root_address : std_logic_vector(13 downto 0);
    signal arrayidx232_674 : std_logic_vector(31 downto 0);
    signal arrayidx255_918 : std_logic_vector(31 downto 0);
    signal arrayidx337_1190 : std_logic_vector(31 downto 0);
    signal arrayidx_467 : std_logic_vector(31 downto 0);
    signal call102_327 : std_logic_vector(7 downto 0);
    signal call106_339 : std_logic_vector(7 downto 0);
    signal call10_74 : std_logic_vector(7 downto 0);
    signal call111_352 : std_logic_vector(7 downto 0);
    signal call115_364 : std_logic_vector(7 downto 0);
    signal call120_377 : std_logic_vector(7 downto 0);
    signal call129_470 : std_logic_vector(7 downto 0);
    signal call133_483 : std_logic_vector(7 downto 0);
    signal call139_501 : std_logic_vector(7 downto 0);
    signal call145_519 : std_logic_vector(7 downto 0);
    signal call14_86 : std_logic_vector(7 downto 0);
    signal call151_537 : std_logic_vector(7 downto 0);
    signal call157_555 : std_logic_vector(7 downto 0);
    signal call163_573 : std_logic_vector(7 downto 0);
    signal call169_591 : std_logic_vector(7 downto 0);
    signal call185_677 : std_logic_vector(7 downto 0);
    signal call189_690 : std_logic_vector(7 downto 0);
    signal call195_708 : std_logic_vector(7 downto 0);
    signal call19_99 : std_logic_vector(7 downto 0);
    signal call201_726 : std_logic_vector(7 downto 0);
    signal call207_744 : std_logic_vector(7 downto 0);
    signal call213_762 : std_logic_vector(7 downto 0);
    signal call219_780 : std_logic_vector(7 downto 0);
    signal call225_798 : std_logic_vector(7 downto 0);
    signal call23_111 : std_logic_vector(7 downto 0);
    signal call261_946 : std_logic_vector(63 downto 0);
    signal call28_124 : std_logic_vector(7 downto 0);
    signal call2_49 : std_logic_vector(7 downto 0);
    signal call312_1099 : std_logic_vector(15 downto 0);
    signal call314_1102 : std_logic_vector(15 downto 0);
    signal call316_1105 : std_logic_vector(15 downto 0);
    signal call318_1108 : std_logic_vector(15 downto 0);
    signal call320_1111 : std_logic_vector(63 downto 0);
    signal call32_136 : std_logic_vector(7 downto 0);
    signal call37_149 : std_logic_vector(7 downto 0);
    signal call41_161 : std_logic_vector(7 downto 0);
    signal call46_174 : std_logic_vector(7 downto 0);
    signal call50_186 : std_logic_vector(7 downto 0);
    signal call55_199 : std_logic_vector(7 downto 0);
    signal call5_61 : std_logic_vector(7 downto 0);
    signal call79_264 : std_logic_vector(7 downto 0);
    signal call84_277 : std_logic_vector(7 downto 0);
    signal call88_289 : std_logic_vector(7 downto 0);
    signal call93_302 : std_logic_vector(7 downto 0);
    signal call97_314 : std_logic_vector(7 downto 0);
    signal call_36 : std_logic_vector(7 downto 0);
    signal cmp180413_408 : std_logic_vector(0 downto 0);
    signal cmp250409_859 : std_logic_vector(0 downto 0);
    signal cmp330406_1131 : std_logic_vector(0 downto 0);
    signal cmp417_393 : std_logic_vector(0 downto 0);
    signal conv100_318 : std_logic_vector(15 downto 0);
    signal conv103_331 : std_logic_vector(15 downto 0);
    signal conv109_343 : std_logic_vector(15 downto 0);
    signal conv112_356 : std_logic_vector(15 downto 0);
    signal conv118_368 : std_logic_vector(15 downto 0);
    signal conv11_78 : std_logic_vector(15 downto 0);
    signal conv121_381 : std_logic_vector(15 downto 0);
    signal conv130_474 : std_logic_vector(63 downto 0);
    signal conv135_487 : std_logic_vector(63 downto 0);
    signal conv141_505 : std_logic_vector(63 downto 0);
    signal conv147_523 : std_logic_vector(63 downto 0);
    signal conv153_541 : std_logic_vector(63 downto 0);
    signal conv159_559 : std_logic_vector(63 downto 0);
    signal conv165_577 : std_logic_vector(63 downto 0);
    signal conv171_595 : std_logic_vector(63 downto 0);
    signal conv17_90 : std_logic_vector(15 downto 0);
    signal conv186_681 : std_logic_vector(63 downto 0);
    signal conv191_694 : std_logic_vector(63 downto 0);
    signal conv197_712 : std_logic_vector(63 downto 0);
    signal conv1_40 : std_logic_vector(15 downto 0);
    signal conv203_730 : std_logic_vector(63 downto 0);
    signal conv209_748 : std_logic_vector(63 downto 0);
    signal conv20_103 : std_logic_vector(15 downto 0);
    signal conv215_766 : std_logic_vector(63 downto 0);
    signal conv221_784 : std_logic_vector(63 downto 0);
    signal conv227_802 : std_logic_vector(63 downto 0);
    signal conv239_835 : std_logic_vector(31 downto 0);
    signal conv241_839 : std_logic_vector(31 downto 0);
    signal conv244_843 : std_logic_vector(31 downto 0);
    signal conv262_952 : std_logic_vector(63 downto 0);
    signal conv26_115 : std_logic_vector(15 downto 0);
    signal conv29_128 : std_logic_vector(15 downto 0);
    signal conv321_1116 : std_logic_vector(63 downto 0);
    signal conv341_1198 : std_logic_vector(7 downto 0);
    signal conv347_1208 : std_logic_vector(7 downto 0);
    signal conv353_1218 : std_logic_vector(7 downto 0);
    signal conv359_1228 : std_logic_vector(7 downto 0);
    signal conv35_140 : std_logic_vector(15 downto 0);
    signal conv365_1238 : std_logic_vector(7 downto 0);
    signal conv371_1248 : std_logic_vector(7 downto 0);
    signal conv377_1258 : std_logic_vector(7 downto 0);
    signal conv383_1268 : std_logic_vector(7 downto 0);
    signal conv38_153 : std_logic_vector(15 downto 0);
    signal conv3_53 : std_logic_vector(15 downto 0);
    signal conv44_165 : std_logic_vector(15 downto 0);
    signal conv47_178 : std_logic_vector(15 downto 0);
    signal conv53_190 : std_logic_vector(15 downto 0);
    signal conv56_203 : std_logic_vector(15 downto 0);
    signal conv61_212 : std_logic_vector(31 downto 0);
    signal conv63_216 : std_logic_vector(31 downto 0);
    signal conv65_220 : std_logic_vector(31 downto 0);
    signal conv69_234 : std_logic_vector(31 downto 0);
    signal conv71_238 : std_logic_vector(31 downto 0);
    signal conv74_242 : std_logic_vector(31 downto 0);
    signal conv77_246 : std_logic_vector(31 downto 0);
    signal conv82_268 : std_logic_vector(15 downto 0);
    signal conv85_281 : std_logic_vector(15 downto 0);
    signal conv8_65 : std_logic_vector(15 downto 0);
    signal conv91_293 : std_logic_vector(15 downto 0);
    signal conv94_306 : std_logic_vector(15 downto 0);
    signal exitcond1_1303 : std_logic_vector(0 downto 0);
    signal exitcond2_822 : std_logic_vector(0 downto 0);
    signal exitcond3_615 : std_logic_vector(0 downto 0);
    signal exitcond_934 : std_logic_vector(0 downto 0);
    signal iNsTr_163_1160 : std_logic_vector(63 downto 0);
    signal iNsTr_25_437 : std_logic_vector(63 downto 0);
    signal iNsTr_38_644 : std_logic_vector(63 downto 0);
    signal iNsTr_52_888 : std_logic_vector(63 downto 0);
    signal indvar429_904 : std_logic_vector(63 downto 0);
    signal indvar443_660 : std_logic_vector(63 downto 0);
    signal indvar459_453 : std_logic_vector(63 downto 0);
    signal indvar_1176 : std_logic_vector(63 downto 0);
    signal indvarx_xnext430_929 : std_logic_vector(63 downto 0);
    signal indvarx_xnext444_817 : std_logic_vector(63 downto 0);
    signal indvarx_xnext460_610 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1298 : std_logic_vector(63 downto 0);
    signal mul242_848 : std_logic_vector(31 downto 0);
    signal mul245_853 : std_logic_vector(31 downto 0);
    signal mul66_230 : std_logic_vector(31 downto 0);
    signal mul72_251 : std_logic_vector(31 downto 0);
    signal mul75_256 : std_logic_vector(31 downto 0);
    signal mul78_261 : std_logic_vector(31 downto 0);
    signal mul_225 : std_logic_vector(31 downto 0);
    signal ptr_deref_1193_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1193_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1193_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1193_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1193_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_602_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_602_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_602_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_602_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_602_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_602_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_809_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_809_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_809_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_809_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_809_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_809_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_920_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_920_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_920_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_920_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_920_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_920_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl101_324 : std_logic_vector(15 downto 0);
    signal shl110_349 : std_logic_vector(15 downto 0);
    signal shl119_374 : std_logic_vector(15 downto 0);
    signal shl132_480 : std_logic_vector(63 downto 0);
    signal shl138_498 : std_logic_vector(63 downto 0);
    signal shl144_516 : std_logic_vector(63 downto 0);
    signal shl150_534 : std_logic_vector(63 downto 0);
    signal shl156_552 : std_logic_vector(63 downto 0);
    signal shl162_570 : std_logic_vector(63 downto 0);
    signal shl168_588 : std_logic_vector(63 downto 0);
    signal shl188_687 : std_logic_vector(63 downto 0);
    signal shl18_96 : std_logic_vector(15 downto 0);
    signal shl194_705 : std_logic_vector(63 downto 0);
    signal shl200_723 : std_logic_vector(63 downto 0);
    signal shl206_741 : std_logic_vector(63 downto 0);
    signal shl212_759 : std_logic_vector(63 downto 0);
    signal shl218_777 : std_logic_vector(63 downto 0);
    signal shl224_795 : std_logic_vector(63 downto 0);
    signal shl27_121 : std_logic_vector(15 downto 0);
    signal shl36_146 : std_logic_vector(15 downto 0);
    signal shl45_171 : std_logic_vector(15 downto 0);
    signal shl54_196 : std_logic_vector(15 downto 0);
    signal shl83_274 : std_logic_vector(15 downto 0);
    signal shl92_299 : std_logic_vector(15 downto 0);
    signal shl9_71 : std_logic_vector(15 downto 0);
    signal shl_46 : std_logic_vector(15 downto 0);
    signal shr344_1204 : std_logic_vector(63 downto 0);
    signal shr350_1214 : std_logic_vector(63 downto 0);
    signal shr356_1224 : std_logic_vector(63 downto 0);
    signal shr362_1234 : std_logic_vector(63 downto 0);
    signal shr368_1244 : std_logic_vector(63 downto 0);
    signal shr374_1254 : std_logic_vector(63 downto 0);
    signal shr380_1264 : std_logic_vector(63 downto 0);
    signal sub_1121 : std_logic_vector(63 downto 0);
    signal tmp338_1194 : std_logic_vector(63 downto 0);
    signal tmp424_1144 : std_logic_vector(31 downto 0);
    signal tmp424x_xop_1156 : std_logic_vector(31 downto 0);
    signal tmp425_1150 : std_logic_vector(0 downto 0);
    signal tmp428_1173 : std_logic_vector(63 downto 0);
    signal tmp436_872 : std_logic_vector(31 downto 0);
    signal tmp436x_xop_884 : std_logic_vector(31 downto 0);
    signal tmp437_878 : std_logic_vector(0 downto 0);
    signal tmp441_901 : std_logic_vector(63 downto 0);
    signal tmp452_628 : std_logic_vector(31 downto 0);
    signal tmp452x_xop_640 : std_logic_vector(31 downto 0);
    signal tmp453_634 : std_logic_vector(0 downto 0);
    signal tmp457_657 : std_logic_vector(63 downto 0);
    signal tmp466_421 : std_logic_vector(31 downto 0);
    signal tmp466x_xop_433 : std_logic_vector(31 downto 0);
    signal tmp467_427 : std_logic_vector(0 downto 0);
    signal tmp471_450 : std_logic_vector(63 downto 0);
    signal type_cast_1114_wire : std_logic_vector(63 downto 0);
    signal type_cast_1129_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1142_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1148_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1154_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1164_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1171_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1179_wire : std_logic_vector(63 downto 0);
    signal type_cast_1182_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1212_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1222_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1232_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1242_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1252_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1262_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1296_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_169_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_194_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_272_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_297_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_322_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_347_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_372_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_390_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_406_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_425_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_431_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_44_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_459_wire : std_logic_vector(63 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_550_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_568_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_586_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_608_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_638_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_655_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_663_wire : std_logic_vector(63 downto 0);
    signal type_cast_666_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_685_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_69_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_703_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_721_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_739_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_793_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_815_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_857_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_876_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_882_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_899_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_910_wire : std_logic_vector(63 downto 0);
    signal type_cast_922_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_927_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_950_wire : std_logic_vector(63 downto 0);
    signal xx_xop473_894 : std_logic_vector(63 downto 0);
    signal xx_xop474_650 : std_logic_vector(63 downto 0);
    signal xx_xop475_443 : std_logic_vector(63 downto 0);
    signal xx_xop_1166 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1188_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1188_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1188_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1188_resized_base_address <= "00000000000000";
    array_obj_ref_465_constant_part_of_offset <= "00000000000000";
    array_obj_ref_465_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_465_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_465_resized_base_address <= "00000000000000";
    array_obj_ref_672_constant_part_of_offset <= "00000100010";
    array_obj_ref_672_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_672_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_672_resized_base_address <= "00000000000";
    array_obj_ref_916_constant_part_of_offset <= "00000000000000";
    array_obj_ref_916_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_916_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_916_resized_base_address <= "00000000000000";
    ptr_deref_1193_word_offset_0 <= "00000000000000";
    ptr_deref_602_word_offset_0 <= "00000000000000";
    ptr_deref_809_word_offset_0 <= "00000000000";
    ptr_deref_920_word_offset_0 <= "00000000000000";
    type_cast_1129_wire_constant <= "00000000000000000000000000000111";
    type_cast_1142_wire_constant <= "00000000000000000000000000000011";
    type_cast_1148_wire_constant <= "00000000000000000000000000000001";
    type_cast_1154_wire_constant <= "11111111111111111111111111111111";
    type_cast_1164_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1171_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1182_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_119_wire_constant <= "0000000000001000";
    type_cast_1202_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1212_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1232_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1242_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1252_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1262_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_144_wire_constant <= "0000000000001000";
    type_cast_169_wire_constant <= "0000000000001000";
    type_cast_194_wire_constant <= "0000000000001000";
    type_cast_272_wire_constant <= "0000000000001000";
    type_cast_297_wire_constant <= "0000000000001000";
    type_cast_322_wire_constant <= "0000000000001000";
    type_cast_347_wire_constant <= "0000000000001000";
    type_cast_372_wire_constant <= "0000000000001000";
    type_cast_390_wire_constant <= "00000000000000000000000000000111";
    type_cast_406_wire_constant <= "00000000000000000000000000000111";
    type_cast_419_wire_constant <= "00000000000000000000000000000011";
    type_cast_425_wire_constant <= "00000000000000000000000000000001";
    type_cast_431_wire_constant <= "11111111111111111111111111111111";
    type_cast_441_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_448_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_44_wire_constant <= "0000000000001000";
    type_cast_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_514_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_550_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_568_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_586_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_608_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_626_wire_constant <= "00000000000000000000000000000011";
    type_cast_632_wire_constant <= "00000000000000000000000000000001";
    type_cast_638_wire_constant <= "11111111111111111111111111111111";
    type_cast_648_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_655_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_666_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_685_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_69_wire_constant <= "0000000000001000";
    type_cast_703_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_721_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_739_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_757_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_775_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_793_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_815_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_857_wire_constant <= "00000000000000000000000000000011";
    type_cast_870_wire_constant <= "00000000000000000000000000000010";
    type_cast_876_wire_constant <= "00000000000000000000000000000001";
    type_cast_882_wire_constant <= "11111111111111111111111111111111";
    type_cast_892_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_899_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_922_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_927_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_94_wire_constant <= "0000000000001000";
    phi_stmt_1176: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1179_wire & type_cast_1182_wire_constant;
      req <= phi_stmt_1176_req_0 & phi_stmt_1176_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1176",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1176_ack_0,
          idata => idata,
          odata => indvar_1176,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1176
    phi_stmt_453: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_457_wire_constant & type_cast_459_wire;
      req <= phi_stmt_453_req_0 & phi_stmt_453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_453",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_453_ack_0,
          idata => idata,
          odata => indvar459_453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_453
    phi_stmt_660: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_663_wire & type_cast_666_wire_constant;
      req <= phi_stmt_660_req_0 & phi_stmt_660_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_660",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_660_ack_0,
          idata => idata,
          odata => indvar443_660,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_660
    phi_stmt_904: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_908_wire_constant & type_cast_910_wire;
      req <= phi_stmt_904_req_0 & phi_stmt_904_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_904",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_904_ack_0,
          idata => idata,
          odata => indvar429_904,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_904
    -- flow-through select operator MUX_1172_inst
    tmp428_1173 <= xx_xop_1166 when (tmp425_1150(0) /=  '0') else type_cast_1171_wire_constant;
    -- flow-through select operator MUX_449_inst
    tmp471_450 <= xx_xop475_443 when (tmp467_427(0) /=  '0') else type_cast_448_wire_constant;
    -- flow-through select operator MUX_656_inst
    tmp457_657 <= xx_xop474_650 when (tmp453_634(0) /=  '0') else type_cast_655_wire_constant;
    -- flow-through select operator MUX_900_inst
    tmp441_901 <= xx_xop473_894 when (tmp437_878(0) /=  '0') else type_cast_899_wire_constant;
    addr_of_1189_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1189_final_reg_req_0;
      addr_of_1189_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1189_final_reg_req_1;
      addr_of_1189_final_reg_ack_1<= rack(0);
      addr_of_1189_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1189_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1188_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx337_1190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_466_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_466_final_reg_req_0;
      addr_of_466_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_466_final_reg_req_1;
      addr_of_466_final_reg_ack_1<= rack(0);
      addr_of_466_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_466_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_465_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_673_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_673_final_reg_req_0;
      addr_of_673_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_673_final_reg_req_1;
      addr_of_673_final_reg_ack_1<= rack(0);
      addr_of_673_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_673_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_672_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx232_674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_917_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_917_final_reg_req_0;
      addr_of_917_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_917_final_reg_req_1;
      addr_of_917_final_reg_ack_1<= rack(0);
      addr_of_917_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_917_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_916_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx255_918,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_102_inst_req_0;
      type_cast_102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_102_inst_req_1;
      type_cast_102_inst_ack_1<= rack(0);
      type_cast_102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1115_inst_req_0;
      type_cast_1115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1115_inst_req_1;
      type_cast_1115_inst_ack_1<= rack(0);
      type_cast_1115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1114_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv321_1116,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_114_inst_req_0;
      type_cast_114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_114_inst_req_1;
      type_cast_114_inst_ack_1<= rack(0);
      type_cast_114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1159_inst_req_0;
      type_cast_1159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1159_inst_req_1;
      type_cast_1159_inst_ack_1<= rack(0);
      type_cast_1159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp424x_xop_1156,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_163_1160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1179_inst_req_0;
      type_cast_1179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1179_inst_req_1;
      type_cast_1179_inst_ack_1<= rack(0);
      type_cast_1179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1179_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1197_inst_req_0;
      type_cast_1197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1197_inst_req_1;
      type_cast_1197_inst_ack_1<= rack(0);
      type_cast_1197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp338_1194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1207_inst_req_0;
      type_cast_1207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1207_inst_req_1;
      type_cast_1207_inst_ack_1<= rack(0);
      type_cast_1207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_1204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_1208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1217_inst_req_0;
      type_cast_1217_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1217_inst_req_1;
      type_cast_1217_inst_ack_1<= rack(0);
      type_cast_1217_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1217_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr350_1214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv353_1218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1227_inst_req_0;
      type_cast_1227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1227_inst_req_1;
      type_cast_1227_inst_ack_1<= rack(0);
      type_cast_1227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr356_1224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv359_1228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1237_inst_req_0;
      type_cast_1237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1237_inst_req_1;
      type_cast_1237_inst_ack_1<= rack(0);
      type_cast_1237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr362_1234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv365_1238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1247_inst_req_0;
      type_cast_1247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1247_inst_req_1;
      type_cast_1247_inst_ack_1<= rack(0);
      type_cast_1247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr368_1244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv371_1248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1257_inst_req_0;
      type_cast_1257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1257_inst_req_1;
      type_cast_1257_inst_ack_1<= rack(0);
      type_cast_1257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr374_1254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv377_1258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1267_inst_req_0;
      type_cast_1267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1267_inst_req_1;
      type_cast_1267_inst_ack_1<= rack(0);
      type_cast_1267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr380_1264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv383_1268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_127_inst_req_0;
      type_cast_127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_127_inst_req_1;
      type_cast_127_inst_ack_1<= rack(0);
      type_cast_127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_152_inst_req_0;
      type_cast_152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_152_inst_req_1;
      type_cast_152_inst_ack_1<= rack(0);
      type_cast_152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_177_inst_req_0;
      type_cast_177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_177_inst_req_1;
      type_cast_177_inst_ack_1<= rack(0);
      type_cast_177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_189_inst_req_0;
      type_cast_189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_189_inst_req_1;
      type_cast_189_inst_ack_1<= rack(0);
      type_cast_189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_202_inst_req_0;
      type_cast_202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_202_inst_req_1;
      type_cast_202_inst_ack_1<= rack(0);
      type_cast_202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_58,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_215_inst_req_0;
      type_cast_215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_215_inst_req_1;
      type_cast_215_inst_ack_1<= rack(0);
      type_cast_215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_83,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_233_inst_req_0;
      type_cast_233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_233_inst_req_1;
      type_cast_233_inst_ack_1<= rack(0);
      type_cast_233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_237_inst_req_0;
      type_cast_237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_237_inst_req_1;
      type_cast_237_inst_ack_1<= rack(0);
      type_cast_237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_241_inst_req_0;
      type_cast_241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_241_inst_req_1;
      type_cast_241_inst_ack_1<= rack(0);
      type_cast_241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_245_inst_req_0;
      type_cast_245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_245_inst_req_1;
      type_cast_245_inst_ack_1<= rack(0);
      type_cast_245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv77_246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_280_inst_req_0;
      type_cast_280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_280_inst_req_1;
      type_cast_280_inst_ack_1<= rack(0);
      type_cast_280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_292_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_292_inst_req_0;
      type_cast_292_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_292_inst_req_1;
      type_cast_292_inst_ack_1<= rack(0);
      type_cast_292_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_292_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_293,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_305_inst_req_0;
      type_cast_305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_305_inst_req_1;
      type_cast_305_inst_ack_1<= rack(0);
      type_cast_305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_317_inst_req_0;
      type_cast_317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_317_inst_req_1;
      type_cast_317_inst_ack_1<= rack(0);
      type_cast_317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_314,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_318,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_330_inst_req_0;
      type_cast_330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_330_inst_req_1;
      type_cast_330_inst_ack_1<= rack(0);
      type_cast_330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call102_327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_342_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_342_inst_req_0;
      type_cast_342_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_342_inst_req_1;
      type_cast_342_inst_ack_1<= rack(0);
      type_cast_342_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_342_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_343,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_355_inst_req_0;
      type_cast_355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_355_inst_req_1;
      type_cast_355_inst_ack_1<= rack(0);
      type_cast_355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_367_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_367_inst_req_0;
      type_cast_367_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_367_inst_req_1;
      type_cast_367_inst_ack_1<= rack(0);
      type_cast_367_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_367_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_380_inst_req_0;
      type_cast_380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_380_inst_req_1;
      type_cast_380_inst_ack_1<= rack(0);
      type_cast_380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call120_377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_39_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_39_inst_req_0;
      type_cast_39_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_39_inst_req_1;
      type_cast_39_inst_ack_1<= rack(0);
      type_cast_39_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_39_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_40,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_436_inst_req_0;
      type_cast_436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_436_inst_req_1;
      type_cast_436_inst_ack_1<= rack(0);
      type_cast_436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp466x_xop_433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_25_437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_459_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_459_inst_req_0;
      type_cast_459_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_459_inst_req_1;
      type_cast_459_inst_ack_1<= rack(0);
      type_cast_459_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_459_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext460_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_459_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_473_inst_req_0;
      type_cast_473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_473_inst_req_1;
      type_cast_473_inst_ack_1<= rack(0);
      type_cast_473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_486_inst_req_0;
      type_cast_486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_486_inst_req_1;
      type_cast_486_inst_ack_1<= rack(0);
      type_cast_486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_504_inst_req_0;
      type_cast_504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_504_inst_req_1;
      type_cast_504_inst_ack_1<= rack(0);
      type_cast_504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_522_inst_req_0;
      type_cast_522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_522_inst_req_1;
      type_cast_522_inst_ack_1<= rack(0);
      type_cast_522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_519,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_52_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_52_inst_req_0;
      type_cast_52_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_52_inst_req_1;
      type_cast_52_inst_ack_1<= rack(0);
      type_cast_52_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_52_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_49,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_540_inst_req_0;
      type_cast_540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_540_inst_req_1;
      type_cast_540_inst_ack_1<= rack(0);
      type_cast_540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_541,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_558_inst_req_0;
      type_cast_558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_558_inst_req_1;
      type_cast_558_inst_ack_1<= rack(0);
      type_cast_558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_559,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_576_inst_req_0;
      type_cast_576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_576_inst_req_1;
      type_cast_576_inst_ack_1<= rack(0);
      type_cast_576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_573,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_594_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_594_inst_req_0;
      type_cast_594_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_594_inst_req_1;
      type_cast_594_inst_ack_1<= rack(0);
      type_cast_594_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_594_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_591,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_595,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp452x_xop_640,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_38_644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_61,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_65,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_663_inst_req_0;
      type_cast_663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_663_inst_req_1;
      type_cast_663_inst_ack_1<= rack(0);
      type_cast_663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext444_817,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_663_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_680_inst_req_0;
      type_cast_680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_680_inst_req_1;
      type_cast_680_inst_ack_1<= rack(0);
      type_cast_680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_680_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call185_677,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_693_inst_req_0;
      type_cast_693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_693_inst_req_1;
      type_cast_693_inst_ack_1<= rack(0);
      type_cast_693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call189_690,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_711_inst_req_0;
      type_cast_711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_711_inst_req_1;
      type_cast_711_inst_ack_1<= rack(0);
      type_cast_711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call195_708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv197_712,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_729_inst_req_0;
      type_cast_729_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_729_inst_req_1;
      type_cast_729_inst_ack_1<= rack(0);
      type_cast_729_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_729_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call201_726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv203_730,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_747_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_747_inst_req_0;
      type_cast_747_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_747_inst_req_1;
      type_cast_747_inst_ack_1<= rack(0);
      type_cast_747_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_747_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call207_744,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv209_748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_765_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_765_inst_req_0;
      type_cast_765_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_765_inst_req_1;
      type_cast_765_inst_ack_1<= rack(0);
      type_cast_765_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_765_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call213_762,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv215_766,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_77_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_77_inst_req_0;
      type_cast_77_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_77_inst_req_1;
      type_cast_77_inst_ack_1<= rack(0);
      type_cast_77_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_77_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_74,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_78,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_783_inst_req_0;
      type_cast_783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_783_inst_req_1;
      type_cast_783_inst_ack_1<= rack(0);
      type_cast_783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call219_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv221_784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_801_inst_req_0;
      type_cast_801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_801_inst_req_1;
      type_cast_801_inst_ack_1<= rack(0);
      type_cast_801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call225_798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv227_802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_834_inst_req_0;
      type_cast_834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_834_inst_req_1;
      type_cast_834_inst_ack_1<= rack(0);
      type_cast_834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv239_835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_838_inst_req_0;
      type_cast_838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_838_inst_req_1;
      type_cast_838_inst_ack_1<= rack(0);
      type_cast_838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add113_361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add122_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv244_843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp436x_xop_884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_89_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_89_inst_req_0;
      type_cast_89_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_89_inst_req_1;
      type_cast_89_inst_ack_1<= rack(0);
      type_cast_89_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_89_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_90,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_910_inst_req_0;
      type_cast_910_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_910_inst_req_1;
      type_cast_910_inst_ack_1<= rack(0);
      type_cast_910_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_910_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext430_929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_910_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_951_inst_req_0;
      type_cast_951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_951_inst_req_1;
      type_cast_951_inst_ack_1<= rack(0);
      type_cast_951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_950_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv262_952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1188_index_1_rename
    process(R_indvar_1187_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1187_resized;
      ov(13 downto 0) := iv;
      R_indvar_1187_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_index_1_resize
    process(indvar_1176) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1176;
      ov := iv(13 downto 0);
      R_indvar_1187_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_root_address_inst
    process(array_obj_ref_1188_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1188_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1188_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_465_index_1_rename
    process(R_indvar459_464_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar459_464_resized;
      ov(13 downto 0) := iv;
      R_indvar459_464_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_465_index_1_resize
    process(indvar459_453) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar459_453;
      ov := iv(13 downto 0);
      R_indvar459_464_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_465_root_address_inst
    process(array_obj_ref_465_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_465_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_465_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_672_index_1_rename
    process(R_indvar443_671_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar443_671_resized;
      ov(10 downto 0) := iv;
      R_indvar443_671_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_672_index_1_resize
    process(indvar443_660) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar443_660;
      ov := iv(10 downto 0);
      R_indvar443_671_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_672_root_address_inst
    process(array_obj_ref_672_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_672_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_672_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_916_index_1_rename
    process(R_indvar429_915_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar429_915_resized;
      ov(13 downto 0) := iv;
      R_indvar429_915_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_916_index_1_resize
    process(indvar429_904) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar429_904;
      ov := iv(13 downto 0);
      R_indvar429_915_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_916_root_address_inst
    process(array_obj_ref_916_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_916_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_916_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1193_addr_0
    process(ptr_deref_1193_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1193_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1193_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1193_base_resize
    process(arrayidx337_1190) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx337_1190;
      ov := iv(13 downto 0);
      ptr_deref_1193_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1193_gather_scatter
    process(ptr_deref_1193_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1193_data_0;
      ov(63 downto 0) := iv;
      tmp338_1194 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1193_root_address_inst
    process(ptr_deref_1193_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1193_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1193_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_addr_0
    process(ptr_deref_602_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_602_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_602_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_base_resize
    process(arrayidx_467) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_467;
      ov := iv(13 downto 0);
      ptr_deref_602_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_gather_scatter
    process(add172_600) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_600;
      ov(63 downto 0) := iv;
      ptr_deref_602_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_602_root_address_inst
    process(ptr_deref_602_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_602_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_602_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_addr_0
    process(ptr_deref_809_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_809_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_809_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_base_resize
    process(arrayidx232_674) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx232_674;
      ov := iv(10 downto 0);
      ptr_deref_809_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_gather_scatter
    process(add228_807) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add228_807;
      ov(63 downto 0) := iv;
      ptr_deref_809_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_809_root_address_inst
    process(ptr_deref_809_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_809_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_809_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_addr_0
    process(ptr_deref_920_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_920_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_920_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_base_resize
    process(arrayidx255_918) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx255_918;
      ov := iv(13 downto 0);
      ptr_deref_920_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_gather_scatter
    process(type_cast_922_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_922_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_920_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_920_root_address_inst
    process(ptr_deref_920_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_920_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_920_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1132_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp330406_1131;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1132_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1132_branch_req_0,
          ack0 => if_stmt_1132_branch_ack_0,
          ack1 => if_stmt_1132_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1304_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1303;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1304_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1304_branch_req_0,
          ack0 => if_stmt_1304_branch_ack_0,
          ack1 => if_stmt_1304_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_394_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp417_393;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_394_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_394_branch_req_0,
          ack0 => if_stmt_394_branch_ack_0,
          ack1 => if_stmt_394_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_409_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp180413_408;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_409_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_409_branch_req_0,
          ack0 => if_stmt_409_branch_ack_0,
          ack1 => if_stmt_409_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_616_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_615;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_616_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_616_branch_req_0,
          ack0 => if_stmt_616_branch_ack_0,
          ack1 => if_stmt_616_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_823_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_822;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_823_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_823_branch_req_0,
          ack0 => if_stmt_823_branch_ack_0,
          ack1 => if_stmt_823_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_860_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp250409_859;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_860_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_860_branch_req_0,
          ack0 => if_stmt_860_branch_ack_0,
          ack1 => if_stmt_860_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_935_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_934;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_935_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_935_branch_req_0,
          ack0 => if_stmt_935_branch_ack_0,
          ack1 => if_stmt_935_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1155_inst
    process(tmp424_1144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp424_1144, type_cast_1154_wire_constant, tmp_var);
      tmp424x_xop_1156 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_432_inst
    process(tmp466_421) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp466_421, type_cast_431_wire_constant, tmp_var);
      tmp466x_xop_433 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_639_inst
    process(tmp452_628) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp452_628, type_cast_638_wire_constant, tmp_var);
      tmp452x_xop_640 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_883_inst
    process(tmp436_872) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp436_872, type_cast_882_wire_constant, tmp_var);
      tmp436x_xop_884 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1165_inst
    process(iNsTr_163_1160) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_163_1160, type_cast_1164_wire_constant, tmp_var);
      xx_xop_1166 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1297_inst
    process(indvar_1176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1176, type_cast_1296_wire_constant, tmp_var);
      indvarx_xnext_1298 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_442_inst
    process(iNsTr_25_437) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_25_437, type_cast_441_wire_constant, tmp_var);
      xx_xop475_443 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_609_inst
    process(indvar459_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar459_453, type_cast_608_wire_constant, tmp_var);
      indvarx_xnext460_610 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_649_inst
    process(iNsTr_38_644) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_38_644, type_cast_648_wire_constant, tmp_var);
      xx_xop474_650 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_816_inst
    process(indvar443_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar443_660, type_cast_815_wire_constant, tmp_var);
      indvarx_xnext444_817 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_893_inst
    process(iNsTr_52_888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_52_888, type_cast_892_wire_constant, tmp_var);
      xx_xop473_894 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_928_inst
    process(indvar429_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar429_904, type_cast_927_wire_constant, tmp_var);
      indvarx_xnext430_929 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1302_inst
    process(indvarx_xnext_1298, tmp428_1173) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1298, tmp428_1173, tmp_var);
      exitcond1_1303 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_614_inst
    process(indvarx_xnext460_610, tmp471_450) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext460_610, tmp471_450, tmp_var);
      exitcond3_615 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_821_inst
    process(indvarx_xnext444_817, tmp457_657) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext444_817, tmp457_657, tmp_var);
      exitcond2_822 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_933_inst
    process(indvarx_xnext430_929, tmp441_901) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext430_929, tmp441_901, tmp_var);
      exitcond_934 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1143_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul245_853, type_cast_1142_wire_constant, tmp_var);
      tmp424_1144 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_420_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_230, type_cast_419_wire_constant, tmp_var);
      tmp466_421 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_627_inst
    process(mul78_261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul78_261, type_cast_626_wire_constant, tmp_var);
      tmp452_628 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_871_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul245_853, type_cast_870_wire_constant, tmp_var);
      tmp436_872 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1203_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1202_wire_constant, tmp_var);
      shr344_1204 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1213_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1212_wire_constant, tmp_var);
      shr350_1214 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1223_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1222_wire_constant, tmp_var);
      shr356_1224 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1233_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1232_wire_constant, tmp_var);
      shr362_1234 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1243_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1242_wire_constant, tmp_var);
      shr368_1244 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1253_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1252_wire_constant, tmp_var);
      shr374_1254 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1263_inst
    process(tmp338_1194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp338_1194, type_cast_1262_wire_constant, tmp_var);
      shr380_1264 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_224_inst
    process(conv63_216, conv61_212) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_216, conv61_212, tmp_var);
      mul_225 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(mul_225, conv65_220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_225, conv65_220, tmp_var);
      mul66_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_250_inst
    process(conv71_238, conv69_234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_238, conv69_234, tmp_var);
      mul72_251 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_255_inst
    process(mul72_251, conv74_242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul72_251, conv74_242, tmp_var);
      mul75_256 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_260_inst
    process(mul75_256, conv77_246) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul75_256, conv77_246, tmp_var);
      mul78_261 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_847_inst
    process(conv241_839, conv239_835) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv241_839, conv239_835, tmp_var);
      mul242_848 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_852_inst
    process(mul242_848, conv244_843) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul242_848, conv244_843, tmp_var);
      mul245_853 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_107_inst
    process(shl18_96, conv20_103) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_96, conv20_103, tmp_var);
      add21_108 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_132_inst
    process(shl27_121, conv29_128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_121, conv29_128, tmp_var);
      add30_133 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_157_inst
    process(shl36_146, conv38_153) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_146, conv38_153, tmp_var);
      add39_158 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_182_inst
    process(shl45_171, conv47_178) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_171, conv47_178, tmp_var);
      add48_183 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_207_inst
    process(shl54_196, conv56_203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_196, conv56_203, tmp_var);
      add57_208 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_285_inst
    process(shl83_274, conv85_281) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_274, conv85_281, tmp_var);
      add86_286 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_310_inst
    process(shl92_299, conv94_306) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_299, conv94_306, tmp_var);
      add95_311 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_335_inst
    process(shl101_324, conv103_331) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl101_324, conv103_331, tmp_var);
      add104_336 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_360_inst
    process(shl110_349, conv112_356) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_349, conv112_356, tmp_var);
      add113_361 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_385_inst
    process(shl119_374, conv121_381) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl119_374, conv121_381, tmp_var);
      add122_386 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_57_inst
    process(shl_46, conv3_53) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_46, conv3_53, tmp_var);
      add_58 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_82_inst
    process(shl9_71, conv11_78) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_71, conv11_78, tmp_var);
      add12_83 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_491_inst
    process(shl132_480, conv135_487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_480, conv135_487, tmp_var);
      add136_492 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_509_inst
    process(shl138_498, conv141_505) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_498, conv141_505, tmp_var);
      add142_510 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_527_inst
    process(shl144_516, conv147_523) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_516, conv147_523, tmp_var);
      add148_528 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_545_inst
    process(shl150_534, conv153_541) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_534, conv153_541, tmp_var);
      add154_546 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_563_inst
    process(shl156_552, conv159_559) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_552, conv159_559, tmp_var);
      add160_564 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_581_inst
    process(shl162_570, conv165_577) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_570, conv165_577, tmp_var);
      add166_582 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_599_inst
    process(shl168_588, conv171_595) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_588, conv171_595, tmp_var);
      add172_600 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_698_inst
    process(shl188_687, conv191_694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl188_687, conv191_694, tmp_var);
      add192_699 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_716_inst
    process(shl194_705, conv197_712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl194_705, conv197_712, tmp_var);
      add198_717 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_734_inst
    process(shl200_723, conv203_730) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl200_723, conv203_730, tmp_var);
      add204_735 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_752_inst
    process(shl206_741, conv209_748) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl206_741, conv209_748, tmp_var);
      add210_753 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_770_inst
    process(shl212_759, conv215_766) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl212_759, conv215_766, tmp_var);
      add216_771 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_788_inst
    process(shl218_777, conv221_784) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl218_777, conv221_784, tmp_var);
      add222_789 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_806_inst
    process(shl224_795, conv227_802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl224_795, conv227_802, tmp_var);
      add228_807 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_120_inst
    process(conv26_115) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_115, type_cast_119_wire_constant, tmp_var);
      shl27_121 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_145_inst
    process(conv35_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_140, type_cast_144_wire_constant, tmp_var);
      shl36_146 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_170_inst
    process(conv44_165) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_165, type_cast_169_wire_constant, tmp_var);
      shl45_171 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_195_inst
    process(conv53_190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_190, type_cast_194_wire_constant, tmp_var);
      shl54_196 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_273_inst
    process(conv82_268) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_268, type_cast_272_wire_constant, tmp_var);
      shl83_274 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_298_inst
    process(conv91_293) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_293, type_cast_297_wire_constant, tmp_var);
      shl92_299 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_323_inst
    process(conv100_318) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv100_318, type_cast_322_wire_constant, tmp_var);
      shl101_324 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_348_inst
    process(conv109_343) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv109_343, type_cast_347_wire_constant, tmp_var);
      shl110_349 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_373_inst
    process(conv118_368) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv118_368, type_cast_372_wire_constant, tmp_var);
      shl119_374 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_45_inst
    process(conv1_40) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_40, type_cast_44_wire_constant, tmp_var);
      shl_46 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_70_inst
    process(conv8_65) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_65, type_cast_69_wire_constant, tmp_var);
      shl9_71 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_95_inst
    process(conv17_90) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_90, type_cast_94_wire_constant, tmp_var);
      shl18_96 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_479_inst
    process(conv130_474) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_474, type_cast_478_wire_constant, tmp_var);
      shl132_480 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_497_inst
    process(add136_492) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_492, type_cast_496_wire_constant, tmp_var);
      shl138_498 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_515_inst
    process(add142_510) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_510, type_cast_514_wire_constant, tmp_var);
      shl144_516 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_533_inst
    process(add148_528) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_528, type_cast_532_wire_constant, tmp_var);
      shl150_534 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_551_inst
    process(add154_546) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_546, type_cast_550_wire_constant, tmp_var);
      shl156_552 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_569_inst
    process(add160_564) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_564, type_cast_568_wire_constant, tmp_var);
      shl162_570 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_587_inst
    process(add166_582) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_582, type_cast_586_wire_constant, tmp_var);
      shl168_588 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_686_inst
    process(conv186_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv186_681, type_cast_685_wire_constant, tmp_var);
      shl188_687 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_704_inst
    process(add192_699) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add192_699, type_cast_703_wire_constant, tmp_var);
      shl194_705 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_722_inst
    process(add198_717) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add198_717, type_cast_721_wire_constant, tmp_var);
      shl200_723 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_740_inst
    process(add204_735) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add204_735, type_cast_739_wire_constant, tmp_var);
      shl206_741 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_758_inst
    process(add210_753) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add210_753, type_cast_757_wire_constant, tmp_var);
      shl212_759 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_776_inst
    process(add216_771) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add216_771, type_cast_775_wire_constant, tmp_var);
      shl218_777 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_794_inst
    process(add222_789) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add222_789, type_cast_793_wire_constant, tmp_var);
      shl224_795 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1120_inst
    process(conv321_1116, conv262_952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv321_1116, conv262_952, tmp_var);
      sub_1121 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1130_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul245_853, type_cast_1129_wire_constant, tmp_var);
      cmp330406_1131 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1149_inst
    process(tmp424_1144) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp424_1144, type_cast_1148_wire_constant, tmp_var);
      tmp425_1150 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_391_inst
    process(mul66_230) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_230, type_cast_390_wire_constant, tmp_var);
      cmp417_393 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_407_inst
    process(mul78_261) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul78_261, type_cast_406_wire_constant, tmp_var);
      cmp180413_408 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_426_inst
    process(tmp466_421) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp466_421, type_cast_425_wire_constant, tmp_var);
      tmp467_427 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_633_inst
    process(tmp452_628) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp452_628, type_cast_632_wire_constant, tmp_var);
      tmp453_634 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_858_inst
    process(mul245_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul245_853, type_cast_857_wire_constant, tmp_var);
      cmp250409_859 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_877_inst
    process(tmp436_872) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp436_872, type_cast_876_wire_constant, tmp_var);
      tmp437_878 <= tmp_var; --
    end process;
    -- shared split operator group (95) : array_obj_ref_1188_index_offset 
    ApIntAdd_group_95: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1187_scaled;
      array_obj_ref_1188_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1188_index_offset_req_0;
      array_obj_ref_1188_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1188_index_offset_req_1;
      array_obj_ref_1188_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_95_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_95_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_95",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 95
    -- shared split operator group (96) : array_obj_ref_465_index_offset 
    ApIntAdd_group_96: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar459_464_scaled;
      array_obj_ref_465_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_465_index_offset_req_0;
      array_obj_ref_465_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_465_index_offset_req_1;
      array_obj_ref_465_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_96_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_96_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : array_obj_ref_672_index_offset 
    ApIntAdd_group_97: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar443_671_scaled;
      array_obj_ref_672_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_672_index_offset_req_0;
      array_obj_ref_672_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_672_index_offset_req_1;
      array_obj_ref_672_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_97_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_97_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- shared split operator group (98) : array_obj_ref_916_index_offset 
    ApIntAdd_group_98: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar429_915_scaled;
      array_obj_ref_916_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_916_index_offset_req_0;
      array_obj_ref_916_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_916_index_offset_req_1;
      array_obj_ref_916_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_98_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_98_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_98",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 98
    -- unary operator type_cast_1114_inst
    process(call320_1111) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call320_1111, tmp_var);
      type_cast_1114_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_950_inst
    process(call261_946) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call261_946, tmp_var);
      type_cast_950_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1193_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1193_load_0_req_0;
      ptr_deref_1193_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1193_load_0_req_1;
      ptr_deref_1193_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1193_word_address_0;
      ptr_deref_1193_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_602_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_602_store_0_req_0;
      ptr_deref_602_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_602_store_0_req_1;
      ptr_deref_602_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_602_word_address_0;
      data_in <= ptr_deref_602_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_809_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_809_store_0_req_0;
      ptr_deref_809_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_809_store_0_req_1;
      ptr_deref_809_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_809_word_address_0;
      data_in <= ptr_deref_809_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_920_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_920_store_0_req_0;
      ptr_deref_920_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_920_store_0_req_1;
      ptr_deref_920_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_920_word_address_0;
      data_in <= ptr_deref_920_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1098_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1098_inst_req_0;
      RPIPE_Block0_done_1098_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1098_inst_req_1;
      RPIPE_Block0_done_1098_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call312_1099 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1101_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1101_inst_req_0;
      RPIPE_Block1_done_1101_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1101_inst_req_1;
      RPIPE_Block1_done_1101_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call314_1102 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1104_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1104_inst_req_0;
      RPIPE_Block2_done_1104_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1104_inst_req_1;
      RPIPE_Block2_done_1104_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call316_1105 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1107_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1107_inst_req_0;
      RPIPE_Block3_done_1107_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1107_inst_req_1;
      RPIPE_Block3_done_1107_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call318_1108 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_288_inst RPIPE_ConvTranspose_input_pipe_123_inst RPIPE_ConvTranspose_input_pipe_160_inst RPIPE_ConvTranspose_input_pipe_198_inst RPIPE_ConvTranspose_input_pipe_148_inst RPIPE_ConvTranspose_input_pipe_98_inst RPIPE_ConvTranspose_input_pipe_313_inst RPIPE_ConvTranspose_input_pipe_48_inst RPIPE_ConvTranspose_input_pipe_185_inst RPIPE_ConvTranspose_input_pipe_110_inst RPIPE_ConvTranspose_input_pipe_85_inst RPIPE_ConvTranspose_input_pipe_173_inst RPIPE_ConvTranspose_input_pipe_263_inst RPIPE_ConvTranspose_input_pipe_73_inst RPIPE_ConvTranspose_input_pipe_35_inst RPIPE_ConvTranspose_input_pipe_135_inst RPIPE_ConvTranspose_input_pipe_301_inst RPIPE_ConvTranspose_input_pipe_276_inst RPIPE_ConvTranspose_input_pipe_676_inst RPIPE_ConvTranspose_input_pipe_725_inst RPIPE_ConvTranspose_input_pipe_707_inst RPIPE_ConvTranspose_input_pipe_743_inst RPIPE_ConvTranspose_input_pipe_689_inst RPIPE_ConvTranspose_input_pipe_590_inst RPIPE_ConvTranspose_input_pipe_572_inst RPIPE_ConvTranspose_input_pipe_554_inst RPIPE_ConvTranspose_input_pipe_536_inst RPIPE_ConvTranspose_input_pipe_518_inst RPIPE_ConvTranspose_input_pipe_500_inst RPIPE_ConvTranspose_input_pipe_482_inst RPIPE_ConvTranspose_input_pipe_469_inst RPIPE_ConvTranspose_input_pipe_338_inst RPIPE_ConvTranspose_input_pipe_60_inst RPIPE_ConvTranspose_input_pipe_326_inst RPIPE_ConvTranspose_input_pipe_376_inst RPIPE_ConvTranspose_input_pipe_363_inst RPIPE_ConvTranspose_input_pipe_351_inst RPIPE_ConvTranspose_input_pipe_761_inst RPIPE_ConvTranspose_input_pipe_779_inst RPIPE_ConvTranspose_input_pipe_797_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_288_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_313_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_263_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_301_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_276_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_676_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_725_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_707_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_743_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_689_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_590_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_572_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_554_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_536_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_518_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_500_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_482_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_469_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_338_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_326_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_376_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_363_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_351_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_761_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_779_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_797_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_288_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_313_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_263_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_301_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_276_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_676_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_725_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_707_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_743_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_689_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_590_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_572_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_554_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_536_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_518_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_500_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_482_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_469_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_338_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_326_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_376_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_363_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_351_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_761_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_779_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_797_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_288_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_160_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_198_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_148_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_98_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_313_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_48_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_185_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_110_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_85_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_173_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_263_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_73_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_35_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_135_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_301_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_276_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_676_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_725_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_707_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_743_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_689_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_590_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_572_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_554_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_536_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_518_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_500_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_482_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_469_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_338_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_60_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_326_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_376_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_363_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_351_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_761_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_779_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_797_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_288_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_160_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_198_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_148_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_98_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_313_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_48_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_185_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_110_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_85_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_173_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_263_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_73_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_35_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_135_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_301_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_276_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_676_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_725_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_707_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_743_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_689_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_590_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_572_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_554_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_536_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_518_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_500_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_482_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_469_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_338_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_60_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_326_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_376_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_363_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_351_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_761_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_779_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_797_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call88_289 <= data_out(319 downto 312);
      call28_124 <= data_out(311 downto 304);
      call41_161 <= data_out(303 downto 296);
      call55_199 <= data_out(295 downto 288);
      call37_149 <= data_out(287 downto 280);
      call19_99 <= data_out(279 downto 272);
      call97_314 <= data_out(271 downto 264);
      call2_49 <= data_out(263 downto 256);
      call50_186 <= data_out(255 downto 248);
      call23_111 <= data_out(247 downto 240);
      call14_86 <= data_out(239 downto 232);
      call46_174 <= data_out(231 downto 224);
      call79_264 <= data_out(223 downto 216);
      call10_74 <= data_out(215 downto 208);
      call_36 <= data_out(207 downto 200);
      call32_136 <= data_out(199 downto 192);
      call93_302 <= data_out(191 downto 184);
      call84_277 <= data_out(183 downto 176);
      call185_677 <= data_out(175 downto 168);
      call201_726 <= data_out(167 downto 160);
      call195_708 <= data_out(159 downto 152);
      call207_744 <= data_out(151 downto 144);
      call189_690 <= data_out(143 downto 136);
      call169_591 <= data_out(135 downto 128);
      call163_573 <= data_out(127 downto 120);
      call157_555 <= data_out(119 downto 112);
      call151_537 <= data_out(111 downto 104);
      call145_519 <= data_out(103 downto 96);
      call139_501 <= data_out(95 downto 88);
      call133_483 <= data_out(87 downto 80);
      call129_470 <= data_out(79 downto 72);
      call106_339 <= data_out(71 downto 64);
      call5_61 <= data_out(63 downto 56);
      call102_327 <= data_out(55 downto 48);
      call120_377 <= data_out(47 downto 40);
      call115_364 <= data_out(39 downto 32);
      call111_352 <= data_out(31 downto 24);
      call213_762 <= data_out(23 downto 16);
      call219_780 <= data_out(15 downto 8);
      call225_798 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_953_inst WPIPE_Block0_start_956_inst WPIPE_Block0_start_959_inst WPIPE_Block0_start_962_inst WPIPE_Block0_start_965_inst WPIPE_Block0_start_968_inst WPIPE_Block0_start_971_inst WPIPE_Block0_start_974_inst WPIPE_Block0_start_977_inst WPIPE_Block0_start_980_inst WPIPE_Block0_start_983_inst WPIPE_Block0_start_986_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block0_start_953_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_956_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_959_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_962_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_965_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_968_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_971_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_974_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_977_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_980_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_983_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_986_inst_req_0;
      WPIPE_Block0_start_953_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_956_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_959_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_962_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_965_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_968_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_971_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_974_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_977_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_980_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_983_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_986_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block0_start_953_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_956_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_959_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_962_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_965_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_968_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_971_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_974_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_977_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_980_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_983_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_986_inst_req_1;
      WPIPE_Block0_start_953_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_956_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_959_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_962_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_965_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_968_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_971_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_974_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_977_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_980_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_983_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_986_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_989_inst WPIPE_Block1_start_992_inst WPIPE_Block1_start_995_inst WPIPE_Block1_start_998_inst WPIPE_Block1_start_1001_inst WPIPE_Block1_start_1004_inst WPIPE_Block1_start_1007_inst WPIPE_Block1_start_1010_inst WPIPE_Block1_start_1013_inst WPIPE_Block1_start_1016_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1022_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block1_start_989_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_992_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_995_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_998_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1001_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1004_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1007_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1010_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1013_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1016_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1022_inst_req_0;
      WPIPE_Block1_start_989_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_992_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_995_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_998_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1001_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1004_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1007_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1010_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1013_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1016_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block1_start_989_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_992_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_995_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_998_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1001_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1004_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1007_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1010_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1013_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1016_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1022_inst_req_1;
      WPIPE_Block1_start_989_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_992_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_995_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_998_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1001_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1004_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1007_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1010_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1013_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1016_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1025_inst WPIPE_Block2_start_1028_inst WPIPE_Block2_start_1031_inst WPIPE_Block2_start_1034_inst WPIPE_Block2_start_1037_inst WPIPE_Block2_start_1040_inst WPIPE_Block2_start_1043_inst WPIPE_Block2_start_1046_inst WPIPE_Block2_start_1049_inst WPIPE_Block2_start_1052_inst WPIPE_Block2_start_1055_inst WPIPE_Block2_start_1058_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block2_start_1025_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1028_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1031_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1034_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1037_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1040_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1043_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1046_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1049_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1052_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1055_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1058_inst_req_0;
      WPIPE_Block2_start_1025_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1028_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1031_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1034_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1037_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1040_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1043_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1046_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1049_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1052_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1055_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1058_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block2_start_1025_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1028_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1031_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1034_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1037_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1040_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1043_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1046_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1049_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1052_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1055_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1058_inst_req_1;
      WPIPE_Block2_start_1025_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1028_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1031_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1034_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1037_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1040_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1043_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1046_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1049_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1052_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1055_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1058_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1061_inst WPIPE_Block3_start_1064_inst WPIPE_Block3_start_1067_inst WPIPE_Block3_start_1070_inst WPIPE_Block3_start_1073_inst WPIPE_Block3_start_1076_inst WPIPE_Block3_start_1079_inst WPIPE_Block3_start_1082_inst WPIPE_Block3_start_1085_inst WPIPE_Block3_start_1088_inst WPIPE_Block3_start_1091_inst WPIPE_Block3_start_1094_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_Block3_start_1061_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1064_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1067_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1070_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1073_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1076_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1079_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1082_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1085_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1088_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1091_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1094_inst_req_0;
      WPIPE_Block3_start_1061_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1064_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1067_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1070_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1073_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1076_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1079_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1082_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1085_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1088_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1091_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1094_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_Block3_start_1061_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1064_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1067_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1070_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1073_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1076_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1079_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1082_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1085_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1088_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1091_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1094_inst_req_1;
      WPIPE_Block3_start_1061_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1064_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1067_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1070_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1073_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1076_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1079_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1082_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1085_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1088_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1091_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1094_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= add_58 & add12_83 & add21_108 & add30_133 & add39_158 & add48_183 & add57_208 & add86_286 & add95_311 & add104_336 & add113_361 & add122_386;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1272_inst WPIPE_ConvTranspose_output_pipe_1284_inst WPIPE_ConvTranspose_output_pipe_1278_inst WPIPE_ConvTranspose_output_pipe_1290_inst WPIPE_ConvTranspose_output_pipe_1287_inst WPIPE_ConvTranspose_output_pipe_1275_inst WPIPE_ConvTranspose_output_pipe_1281_inst WPIPE_ConvTranspose_output_pipe_1269_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1272_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1278_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1275_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1269_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1272_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1278_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1275_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1269_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1272_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1284_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1278_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1275_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1281_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1269_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1272_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1284_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1278_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1275_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1281_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1269_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv377_1258 & conv353_1218 & conv365_1238 & conv341_1198 & conv347_1208 & conv371_1248 & conv359_1228 & conv383_1268;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1122_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1122_inst_req_0;
      WPIPE_elapsed_time_pipe_1122_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1122_inst_req_1;
      WPIPE_elapsed_time_pipe_1122_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1121;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_946_call call_stmt_1111_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_946_call_req_0;
      reqL_unguarded(0) <= call_stmt_1111_call_req_0;
      call_stmt_946_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1111_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_946_call_req_1;
      reqR_unguarded(0) <= call_stmt_1111_call_req_1;
      call_stmt_946_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1111_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call261_946 <= data_out(127 downto 64);
      call320_1111 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3357_start: Boolean;
  signal convTransposeA_CP_3357_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1477_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1320_inst_ack_0 : boolean;
  signal phi_stmt_1471_ack_0 : boolean;
  signal RPIPE_Block0_start_1326_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1335_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_req_0 : boolean;
  signal type_cast_1624_inst_ack_1 : boolean;
  signal type_cast_1477_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1323_inst_ack_1 : boolean;
  signal phi_stmt_1404_req_0 : boolean;
  signal RPIPE_Block0_start_1320_inst_req_1 : boolean;
  signal type_cast_1598_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1320_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1326_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1320_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1338_inst_req_1 : boolean;
  signal phi_stmt_1471_req_1 : boolean;
  signal if_stmt_1631_branch_req_0 : boolean;
  signal RPIPE_Block0_start_1323_inst_req_0 : boolean;
  signal type_cast_1624_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1323_inst_ack_0 : boolean;
  signal phi_stmt_1411_req_0 : boolean;
  signal RPIPE_Block0_start_1326_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1329_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1329_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1323_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1329_inst_req_1 : boolean;
  signal if_stmt_1631_branch_ack_1 : boolean;
  signal RPIPE_Block0_start_1329_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1332_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1332_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1332_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1332_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1335_inst_ack_0 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal type_cast_1477_inst_ack_0 : boolean;
  signal type_cast_1477_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1341_inst_req_1 : boolean;
  signal type_cast_1598_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1341_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1341_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1639_inst_req_1 : boolean;
  signal phi_stmt_1471_req_0 : boolean;
  signal phi_stmt_1411_ack_0 : boolean;
  signal type_cast_1417_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1350_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1350_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1350_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1350_inst_ack_1 : boolean;
  signal type_cast_1598_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1344_inst_req_0 : boolean;
  signal type_cast_1598_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1341_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1338_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1338_inst_ack_0 : boolean;
  signal phi_stmt_1404_ack_0 : boolean;
  signal RPIPE_Block0_start_1326_inst_ack_1 : boolean;
  signal WPIPE_Block0_done_1639_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1338_inst_ack_1 : boolean;
  signal phi_stmt_1411_req_1 : boolean;
  signal RPIPE_Block0_start_1344_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1344_inst_ack_1 : boolean;
  signal type_cast_1624_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1347_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1347_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1639_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1347_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1347_inst_ack_1 : boolean;
  signal type_cast_1417_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1344_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1353_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1353_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1353_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1353_inst_ack_1 : boolean;
  signal type_cast_1624_inst_req_0 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal type_cast_1358_inst_req_0 : boolean;
  signal type_cast_1358_inst_ack_0 : boolean;
  signal type_cast_1358_inst_req_1 : boolean;
  signal type_cast_1358_inst_ack_1 : boolean;
  signal WPIPE_Block0_done_1639_inst_req_0 : boolean;
  signal type_cast_1417_inst_ack_0 : boolean;
  signal type_cast_1362_inst_req_0 : boolean;
  signal type_cast_1362_inst_ack_0 : boolean;
  signal type_cast_1362_inst_req_1 : boolean;
  signal type_cast_1362_inst_ack_1 : boolean;
  signal type_cast_1417_inst_req_0 : boolean;
  signal type_cast_1372_inst_req_0 : boolean;
  signal type_cast_1372_inst_ack_0 : boolean;
  signal type_cast_1372_inst_req_1 : boolean;
  signal type_cast_1372_inst_ack_1 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal type_cast_1499_inst_req_0 : boolean;
  signal type_cast_1499_inst_ack_0 : boolean;
  signal type_cast_1499_inst_req_1 : boolean;
  signal type_cast_1499_inst_ack_1 : boolean;
  signal type_cast_1513_inst_req_0 : boolean;
  signal type_cast_1513_inst_ack_0 : boolean;
  signal type_cast_1513_inst_req_1 : boolean;
  signal type_cast_1513_inst_ack_1 : boolean;
  signal if_stmt_1631_branch_ack_0 : boolean;
  signal phi_stmt_1404_req_1 : boolean;
  signal type_cast_1410_inst_ack_1 : boolean;
  signal type_cast_1410_inst_req_1 : boolean;
  signal type_cast_1410_inst_ack_0 : boolean;
  signal type_cast_1410_inst_req_0 : boolean;
  signal array_obj_ref_1519_index_offset_req_0 : boolean;
  signal array_obj_ref_1519_index_offset_ack_0 : boolean;
  signal array_obj_ref_1519_index_offset_req_1 : boolean;
  signal array_obj_ref_1519_index_offset_ack_1 : boolean;
  signal addr_of_1520_final_reg_req_0 : boolean;
  signal addr_of_1520_final_reg_ack_0 : boolean;
  signal addr_of_1520_final_reg_req_1 : boolean;
  signal addr_of_1520_final_reg_ack_1 : boolean;
  signal ptr_deref_1524_load_0_req_0 : boolean;
  signal ptr_deref_1524_load_0_ack_0 : boolean;
  signal ptr_deref_1524_load_0_req_1 : boolean;
  signal ptr_deref_1524_load_0_ack_1 : boolean;
  signal type_cast_1529_inst_req_0 : boolean;
  signal type_cast_1529_inst_ack_0 : boolean;
  signal type_cast_1529_inst_req_1 : boolean;
  signal type_cast_1529_inst_ack_1 : boolean;
  signal type_cast_1543_inst_req_0 : boolean;
  signal type_cast_1543_inst_ack_0 : boolean;
  signal type_cast_1543_inst_req_1 : boolean;
  signal type_cast_1543_inst_ack_1 : boolean;
  signal array_obj_ref_1549_index_offset_req_0 : boolean;
  signal array_obj_ref_1549_index_offset_ack_0 : boolean;
  signal array_obj_ref_1549_index_offset_req_1 : boolean;
  signal array_obj_ref_1549_index_offset_ack_1 : boolean;
  signal addr_of_1550_final_reg_req_0 : boolean;
  signal addr_of_1550_final_reg_ack_0 : boolean;
  signal addr_of_1550_final_reg_req_1 : boolean;
  signal addr_of_1550_final_reg_ack_1 : boolean;
  signal ptr_deref_1553_store_0_req_0 : boolean;
  signal ptr_deref_1553_store_0_ack_0 : boolean;
  signal ptr_deref_1553_store_0_req_1 : boolean;
  signal ptr_deref_1553_store_0_ack_1 : boolean;
  signal type_cast_1559_inst_req_0 : boolean;
  signal type_cast_1559_inst_ack_0 : boolean;
  signal type_cast_1559_inst_req_1 : boolean;
  signal type_cast_1559_inst_ack_1 : boolean;
  signal if_stmt_1574_branch_req_0 : boolean;
  signal if_stmt_1574_branch_ack_1 : boolean;
  signal if_stmt_1574_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3357_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3357_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3357_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3357_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3357: Block -- control-path 
    signal convTransposeA_CP_3357_elements: BooleanArray(87 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3357_elements(0) <= convTransposeA_CP_3357_start;
    convTransposeA_CP_3357_symbol <= convTransposeA_CP_3357_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354__entry__
      -- CP-element group 0: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1318/branch_block_stmt_1318__entry__
      -- CP-element group 0: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/$entry
      -- CP-element group 0: 	 branch_block_stmt_1318/$entry
      -- 
    rr_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(0), ack => RPIPE_Block0_start_1320_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Update/$entry
      -- 
    ra_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1320_inst_ack_0, ack => convTransposeA_CP_3357_elements(1)); -- 
    cr_3410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(1), ack => RPIPE_Block0_start_1320_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1320_Update/$exit
      -- 
    ca_3411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1320_inst_ack_1, ack => convTransposeA_CP_3357_elements(2)); -- 
    rr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(2), ack => RPIPE_Block0_start_1323_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Update/cr
      -- 
    ra_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1323_inst_ack_0, ack => convTransposeA_CP_3357_elements(3)); -- 
    cr_3424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(3), ack => RPIPE_Block0_start_1323_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1323_Update/ca
      -- 
    ca_3425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1323_inst_ack_1, ack => convTransposeA_CP_3357_elements(4)); -- 
    rr_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(4), ack => RPIPE_Block0_start_1326_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Sample/ra
      -- 
    ra_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1326_inst_ack_0, ack => convTransposeA_CP_3357_elements(5)); -- 
    cr_3438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(5), ack => RPIPE_Block0_start_1326_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1326_Update/ca
      -- 
    ca_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1326_inst_ack_1, ack => convTransposeA_CP_3357_elements(6)); -- 
    rr_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(6), ack => RPIPE_Block0_start_1329_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_update_start_
      -- 
    ra_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1329_inst_ack_0, ack => convTransposeA_CP_3357_elements(7)); -- 
    cr_3452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(7), ack => RPIPE_Block0_start_1329_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1329_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Sample/rr
      -- 
    ca_3453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1329_inst_ack_1, ack => convTransposeA_CP_3357_elements(8)); -- 
    rr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(8), ack => RPIPE_Block0_start_1332_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Update/cr
      -- 
    ra_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1332_inst_ack_0, ack => convTransposeA_CP_3357_elements(9)); -- 
    cr_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(9), ack => RPIPE_Block0_start_1332_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1332_Update/ca
      -- 
    ca_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1332_inst_ack_1, ack => convTransposeA_CP_3357_elements(10)); -- 
    rr_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(10), ack => RPIPE_Block0_start_1335_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Sample/ra
      -- 
    ra_3476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1335_inst_ack_0, ack => convTransposeA_CP_3357_elements(11)); -- 
    cr_3480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(11), ack => RPIPE_Block0_start_1335_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1335_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Sample/$entry
      -- 
    ca_3481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1335_inst_ack_1, ack => convTransposeA_CP_3357_elements(12)); -- 
    rr_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(12), ack => RPIPE_Block0_start_1338_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Sample/$exit
      -- 
    ra_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1338_inst_ack_0, ack => convTransposeA_CP_3357_elements(13)); -- 
    cr_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(13), ack => RPIPE_Block0_start_1338_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1338_Update/ca
      -- 
    ca_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1338_inst_ack_1, ack => convTransposeA_CP_3357_elements(14)); -- 
    rr_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(14), ack => RPIPE_Block0_start_1341_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_update_start_
      -- 
    ra_3504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1341_inst_ack_0, ack => convTransposeA_CP_3357_elements(15)); -- 
    cr_3508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(15), ack => RPIPE_Block0_start_1341_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1341_Update/ca
      -- 
    ca_3509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1341_inst_ack_1, ack => convTransposeA_CP_3357_elements(16)); -- 
    rr_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(16), ack => RPIPE_Block0_start_1344_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Update/$entry
      -- 
    ra_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1344_inst_ack_0, ack => convTransposeA_CP_3357_elements(17)); -- 
    cr_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(17), ack => RPIPE_Block0_start_1344_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1344_Update/$exit
      -- 
    ca_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1344_inst_ack_1, ack => convTransposeA_CP_3357_elements(18)); -- 
    rr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(18), ack => RPIPE_Block0_start_1347_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/cr
      -- 
    ra_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1347_inst_ack_0, ack => convTransposeA_CP_3357_elements(19)); -- 
    cr_3536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(19), ack => RPIPE_Block0_start_1347_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1347_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_sample_start_
      -- 
    ca_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1347_inst_ack_1, ack => convTransposeA_CP_3357_elements(20)); -- 
    rr_3545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(20), ack => RPIPE_Block0_start_1350_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_sample_completed_
      -- 
    ra_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1350_inst_ack_0, ack => convTransposeA_CP_3357_elements(21)); -- 
    cr_3550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(21), ack => RPIPE_Block0_start_1350_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1350_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/rr
      -- 
    ca_3551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1350_inst_ack_1, ack => convTransposeA_CP_3357_elements(22)); -- 
    rr_3559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(22), ack => RPIPE_Block0_start_1353_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/cr
      -- 
    ra_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1353_inst_ack_0, ack => convTransposeA_CP_3357_elements(23)); -- 
    cr_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(23), ack => RPIPE_Block0_start_1353_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/$exit
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354__exit__
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401__entry__
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1321_to_assign_stmt_1354/RPIPE_Block0_start_1353_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Update/cr
      -- 
    ca_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1353_inst_ack_1, ack => convTransposeA_CP_3357_elements(24)); -- 
    rr_3576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(24), ack => type_cast_1358_inst_req_0); -- 
    cr_3581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(24), ack => type_cast_1358_inst_req_1); -- 
    rr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(24), ack => type_cast_1362_inst_req_0); -- 
    cr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(24), ack => type_cast_1362_inst_req_1); -- 
    rr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(24), ack => type_cast_1372_inst_req_0); -- 
    cr_3609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(24), ack => type_cast_1372_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Sample/ra
      -- 
    ra_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_0, ack => convTransposeA_CP_3357_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1358_Update/ca
      -- 
    ca_3582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_1, ack => convTransposeA_CP_3357_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Sample/ra
      -- 
    ra_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1362_inst_ack_0, ack => convTransposeA_CP_3357_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1362_Update/ca
      -- 
    ca_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1362_inst_ack_1, ack => convTransposeA_CP_3357_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Sample/ra
      -- 
    ra_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1372_inst_ack_0, ack => convTransposeA_CP_3357_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/type_cast_1372_Update/ca
      -- 
    ca_3610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1372_inst_ack_1, ack => convTransposeA_CP_3357_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31:  members (8) 
      -- CP-element group 31: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/$entry
      -- CP-element group 31: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/$entry
      -- CP-element group 31: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401__exit__
      -- CP-element group 31: 	 branch_block_stmt_1318/assign_stmt_1359_to_assign_stmt_1401/$exit
      -- 
    convTransposeA_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(26) & convTransposeA_CP_3357_elements(28) & convTransposeA_CP_3357_elements(30);
      gj_convTransposeA_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	87 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Sample/ra
      -- 
    ra_3625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1499_inst_ack_0, ack => convTransposeA_CP_3357_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	87 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Sample/rr
      -- 
    ca_3630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1499_inst_ack_1, ack => convTransposeA_CP_3357_elements(33)); -- 
    rr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(33), ack => type_cast_1513_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Sample/ra
      -- 
    ra_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_0, ack => convTransposeA_CP_3357_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	87 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Sample/req
      -- 
    ca_3644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_1, ack => convTransposeA_CP_3357_elements(35)); -- 
    req_3669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(35), ack => array_obj_ref_1519_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Sample/ack
      -- 
    ack_3670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1519_index_offset_ack_0, ack => convTransposeA_CP_3357_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	87 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_request/req
      -- 
    ack_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1519_index_offset_ack_1, ack => convTransposeA_CP_3357_elements(37)); -- 
    req_3684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(37), ack => addr_of_1520_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_request/ack
      -- 
    ack_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1520_final_reg_ack_0, ack => convTransposeA_CP_3357_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	87 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/word_access_start/word_0/rr
      -- 
    ack_3690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1520_final_reg_ack_1, ack => convTransposeA_CP_3357_elements(39)); -- 
    rr_3723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(39), ack => ptr_deref_1524_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Sample/word_access_start/word_0/ra
      -- 
    ra_3724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1524_load_0_ack_0, ack => convTransposeA_CP_3357_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	87 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/ptr_deref_1524_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/ptr_deref_1524_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/ptr_deref_1524_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/ptr_deref_1524_Merge/merge_ack
      -- 
    ca_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1524_load_0_ack_1, ack => convTransposeA_CP_3357_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	87 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Sample/ra
      -- 
    ra_3749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1529_inst_ack_0, ack => convTransposeA_CP_3357_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	87 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Sample/rr
      -- 
    ca_3754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1529_inst_ack_1, ack => convTransposeA_CP_3357_elements(43)); -- 
    rr_3762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(43), ack => type_cast_1543_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Sample/ra
      -- 
    ra_3763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1543_inst_ack_0, ack => convTransposeA_CP_3357_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	87 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Sample/req
      -- 
    ca_3768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1543_inst_ack_1, ack => convTransposeA_CP_3357_elements(45)); -- 
    req_3793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(45), ack => array_obj_ref_1549_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Sample/ack
      -- 
    ack_3794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1549_index_offset_ack_0, ack => convTransposeA_CP_3357_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	87 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_request/req
      -- 
    ack_3799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1549_index_offset_ack_1, ack => convTransposeA_CP_3357_elements(47)); -- 
    req_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(47), ack => addr_of_1550_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_request/ack
      -- 
    ack_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1550_final_reg_ack_0, ack => convTransposeA_CP_3357_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	87 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_word_addrgen/root_register_ack
      -- 
    ack_3814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1550_final_reg_ack_1, ack => convTransposeA_CP_3357_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	41 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/ptr_deref_1553_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/ptr_deref_1553_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/ptr_deref_1553_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/ptr_deref_1553_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/word_access_start/word_0/rr
      -- 
    rr_3852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(50), ack => ptr_deref_1553_store_0_req_0); -- 
    convTransposeA_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(49) & convTransposeA_CP_3357_elements(41);
      gj_convTransposeA_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Sample/word_access_start/word_0/ra
      -- 
    ra_3853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1553_store_0_ack_0, ack => convTransposeA_CP_3357_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	87 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/word_access_complete/word_0/ca
      -- 
    ca_3864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1553_store_0_ack_1, ack => convTransposeA_CP_3357_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	87 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Sample/ra
      -- 
    ra_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_0, ack => convTransposeA_CP_3357_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	87 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Update/ca
      -- 
    ca_3878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_1, ack => convTransposeA_CP_3357_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	36 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574__entry__
      -- CP-element group 55: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573__exit__
      -- CP-element group 55: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/$exit
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1318/R_cmp_1575_place
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1318/if_stmt_1574_else_link/$entry
      -- 
    branch_req_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(55), ack => if_stmt_1574_branch_req_0); -- 
    convTransposeA_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(46) & convTransposeA_CP_3357_elements(52) & convTransposeA_CP_3357_elements(54) & convTransposeA_CP_3357_elements(36);
      gj_convTransposeA_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	82 
    -- CP-element group 56: 	83 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1318/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/merge_stmt_1580_PhiAck/dummy
      -- CP-element group 56: 	 branch_block_stmt_1318/merge_stmt_1580_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/assign_stmt_1586__entry__
      -- CP-element group 56: 	 branch_block_stmt_1318/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/assign_stmt_1586__exit__
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1318/merge_stmt_1580_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/merge_stmt_1580_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1318/merge_stmt_1580__exit__
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/if_stmt_1574_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1318/if_stmt_1574_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1318/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1318/assign_stmt_1586/$entry
      -- CP-element group 56: 	 branch_block_stmt_1318/assign_stmt_1586/$exit
      -- 
    if_choice_transition_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1574_branch_ack_1, ack => convTransposeA_CP_3357_elements(56)); -- 
    cr_4079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(56), ack => type_cast_1477_inst_req_1); -- 
    rr_4074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(56), ack => type_cast_1477_inst_req_0); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1318/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1318/merge_stmt_1588_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/merge_stmt_1588__exit__
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630__entry__
      -- CP-element group 57: 	 branch_block_stmt_1318/merge_stmt_1588_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1318/merge_stmt_1588_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1318/merge_stmt_1588_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1318/if_stmt_1574_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1318/if_stmt_1574_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1318/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/$entry
      -- CP-element group 57: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_sample_start_
      -- 
    else_choice_transition_3895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1574_branch_ack_0, ack => convTransposeA_CP_3357_elements(57)); -- 
    rr_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(57), ack => type_cast_1598_inst_req_0); -- 
    cr_3916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(57), ack => type_cast_1598_inst_req_1); -- 
    cr_3944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(57), ack => type_cast_1624_inst_req_1); -- 
    cr_3930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(57), ack => type_cast_1607_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_sample_completed_
      -- 
    ra_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_0, ack => convTransposeA_CP_3357_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1598_update_completed_
      -- 
    ca_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_1, ack => convTransposeA_CP_3357_elements(59)); -- 
    rr_3925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(59), ack => type_cast_1607_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Sample/ra
      -- 
    ra_3926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => convTransposeA_CP_3357_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1607_Update/$exit
      -- 
    ca_3931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => convTransposeA_CP_3357_elements(61)); -- 
    rr_3939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(61), ack => type_cast_1624_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_sample_completed_
      -- 
    ra_3940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1624_inst_ack_0, ack => convTransposeA_CP_3357_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631__entry__
      -- CP-element group 63: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630__exit__
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/type_cast_1624_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1318/R_cmp116_1632_place
      -- CP-element group 63: 	 branch_block_stmt_1318/if_stmt_1631_else_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1318/assign_stmt_1594_to_assign_stmt_1630/$exit
      -- 
    ca_3945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1624_inst_ack_1, ack => convTransposeA_CP_3357_elements(63)); -- 
    branch_req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(63), ack => if_stmt_1631_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1318/if_stmt_1631_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1318/merge_stmt_1637__exit__
      -- CP-element group 64: 	 branch_block_stmt_1318/if_stmt_1631_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1318/assign_stmt_1642__entry__
      -- CP-element group 64: 	 branch_block_stmt_1318/merge_stmt_1637_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1318/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1318/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1318/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1318/assign_stmt_1642/$entry
      -- CP-element group 64: 	 branch_block_stmt_1318/merge_stmt_1637_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_1318/merge_stmt_1637_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1318/merge_stmt_1637_PhiAck/$entry
      -- 
    if_choice_transition_3958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1631_branch_ack_1, ack => convTransposeA_CP_3357_elements(64)); -- 
    req_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(64), ack => WPIPE_Block0_done_1639_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	71 
    -- CP-element group 65: 	72 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	75 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/if_stmt_1631_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1318/if_stmt_1631_else_link/$exit
      -- 
    else_choice_transition_3962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1631_branch_ack_0, ack => convTransposeA_CP_3357_elements(65)); -- 
    cr_4047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(65), ack => type_cast_1417_inst_req_1); -- 
    rr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(65), ack => type_cast_1417_inst_req_0); -- 
    cr_4024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(65), ack => type_cast_1410_inst_req_1); -- 
    rr_4019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(65), ack => type_cast_1410_inst_req_0); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Update/req
      -- CP-element group 66: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_sample_completed_
      -- 
    ack_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1639_inst_ack_0, ack => convTransposeA_CP_3357_elements(66)); -- 
    req_3980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(66), ack => WPIPE_Block0_done_1639_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1318/branch_block_stmt_1318__exit__
      -- CP-element group 67: 	 branch_block_stmt_1318/$exit
      -- CP-element group 67: 	 branch_block_stmt_1318/merge_stmt_1644__exit__
      -- CP-element group 67: 	 branch_block_stmt_1318/return__
      -- CP-element group 67: 	 branch_block_stmt_1318/assign_stmt_1642__exit__
      -- CP-element group 67: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1318/merge_stmt_1644_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1318/assign_stmt_1642/WPIPE_Block0_done_1639_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1318/assign_stmt_1642/$exit
      -- CP-element group 67: 	 branch_block_stmt_1318/merge_stmt_1644_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_1318/merge_stmt_1644_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1318/merge_stmt_1644_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1318/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1318/return___PhiReq/$entry
      -- 
    ack_3981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1639_inst_ack_1, ack => convTransposeA_CP_3357_elements(67)); -- 
    -- CP-element group 68:  transition  output  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_req
      -- CP-element group 68: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/$exit
      -- CP-element group 68: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1408_konst_delay_trans
      -- 
    phi_stmt_1404_req_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1404_req_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(68), ack => phi_stmt_1404_req_0); -- 
    -- Element group convTransposeA_CP_3357_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => convTransposeA_CP_3357_elements(31), ack => convTransposeA_CP_3357_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1415_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_req
      -- CP-element group 69: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/$exit
      -- 
    phi_stmt_1411_req_4000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1411_req_4000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(69), ack => phi_stmt_1411_req_0); -- 
    -- Element group convTransposeA_CP_3357_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_3357_elements(31), ack => convTransposeA_CP_3357_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  transition  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1318/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(68) & convTransposeA_CP_3357_elements(69);
      gj_convTransposeA_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	65 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Sample/$exit
      -- 
    ra_4020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1410_inst_ack_0, ack => convTransposeA_CP_3357_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	65 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/Update/$exit
      -- 
    ca_4025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1410_inst_ack_1, ack => convTransposeA_CP_3357_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/$exit
      -- CP-element group 73: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/type_cast_1410/$exit
      -- CP-element group 73: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1404/phi_stmt_1404_req
      -- 
    phi_stmt_1404_req_4026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1404_req_4026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(73), ack => phi_stmt_1404_req_1); -- 
    convTransposeA_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(71) & convTransposeA_CP_3357_elements(72);
      gj_convTransposeA_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Sample/$exit
      -- 
    ra_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_0, ack => convTransposeA_CP_3357_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Update/ca
      -- CP-element group 75: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/Update/$exit
      -- 
    ca_4048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_1, ack => convTransposeA_CP_3357_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_req
      -- CP-element group 76: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/type_cast_1417/$exit
      -- CP-element group 76: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/phi_stmt_1411_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1411/$exit
      -- 
    phi_stmt_1411_req_4049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1411_req_4049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(76), ack => phi_stmt_1411_req_1); -- 
    convTransposeA_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(74) & convTransposeA_CP_3357_elements(75);
      gj_convTransposeA_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1318/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(73) & convTransposeA_CP_3357_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  merge  fork  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1318/merge_stmt_1403_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1318/merge_stmt_1403_PhiReqMerge
      -- 
    convTransposeA_CP_3357_elements(78) <= OrReduce(convTransposeA_CP_3357_elements(70) & convTransposeA_CP_3357_elements(77));
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1318/merge_stmt_1403_PhiAck/phi_stmt_1404_ack
      -- 
    phi_stmt_1404_ack_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1404_ack_0, ack => convTransposeA_CP_3357_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1318/merge_stmt_1403_PhiAck/phi_stmt_1411_ack
      -- 
    phi_stmt_1411_ack_4055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1411_ack_0, ack => convTransposeA_CP_3357_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (10) 
      -- CP-element group 81: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 81: 	 branch_block_stmt_1318/assign_stmt_1423_to_assign_stmt_1468__exit__
      -- CP-element group 81: 	 branch_block_stmt_1318/assign_stmt_1423_to_assign_stmt_1468__entry__
      -- CP-element group 81: 	 branch_block_stmt_1318/merge_stmt_1403__exit__
      -- CP-element group 81: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1471/$entry
      -- CP-element group 81: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$entry
      -- CP-element group 81: 	 branch_block_stmt_1318/merge_stmt_1403_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_1318/assign_stmt_1423_to_assign_stmt_1468/$entry
      -- CP-element group 81: 	 branch_block_stmt_1318/assign_stmt_1423_to_assign_stmt_1468/$exit
      -- 
    convTransposeA_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(79) & convTransposeA_CP_3357_elements(80);
      gj_convTransposeA_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	56 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/ra
      -- 
    ra_4075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1477_inst_ack_0, ack => convTransposeA_CP_3357_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	56 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/ca
      -- CP-element group 83: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/$exit
      -- 
    ca_4080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1477_inst_ack_1, ack => convTransposeA_CP_3357_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_req
      -- CP-element group 84: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/$exit
      -- CP-element group 84: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1471/$exit
      -- CP-element group 84: 	 branch_block_stmt_1318/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1471_req_4081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1471_req_4081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(84), ack => phi_stmt_1471_req_1); -- 
    convTransposeA_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3357_elements(82) & convTransposeA_CP_3357_elements(83);
      gj_convTransposeA_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3357_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  output  delay-element  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1475_konst_delay_trans
      -- CP-element group 85: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1471/$exit
      -- CP-element group 85: 	 branch_block_stmt_1318/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1471/phi_stmt_1471_req
      -- 
    phi_stmt_1471_req_4092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1471_req_4092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(85), ack => phi_stmt_1471_req_0); -- 
    -- Element group convTransposeA_CP_3357_elements(85) is a control-delay.
    cp_element_85_delay: control_delay_element  generic map(name => " 85_delay", delay_value => 1)  port map(req => convTransposeA_CP_3357_elements(81), ack => convTransposeA_CP_3357_elements(85), clk => clk, reset =>reset);
    -- CP-element group 86:  merge  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1318/merge_stmt_1470_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_1318/merge_stmt_1470_PhiAck/$entry
      -- 
    convTransposeA_CP_3357_elements(86) <= OrReduce(convTransposeA_CP_3357_elements(84) & convTransposeA_CP_3357_elements(85));
    -- CP-element group 87:  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	47 
    -- CP-element group 87: 	49 
    -- CP-element group 87: 	52 
    -- CP-element group 87: 	53 
    -- CP-element group 87: 	54 
    -- CP-element group 87: 	32 
    -- CP-element group 87: 	33 
    -- CP-element group 87: 	35 
    -- CP-element group 87: 	37 
    -- CP-element group 87: 	39 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	42 
    -- CP-element group 87: 	43 
    -- CP-element group 87: 	45 
    -- CP-element group 87:  members (51) 
      -- CP-element group 87: 	 branch_block_stmt_1318/merge_stmt_1470_PhiAck/phi_stmt_1471_ack
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573__entry__
      -- CP-element group 87: 	 branch_block_stmt_1318/merge_stmt_1470__exit__
      -- CP-element group 87: 	 branch_block_stmt_1318/merge_stmt_1470_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1499_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1513_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1519_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1520_complete/req
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1524_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1529_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1543_Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_update_start
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/array_obj_ref_1549_final_index_sum_regn_Update/req
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/addr_of_1550_complete/req
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/word_access_complete/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/word_access_complete/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/ptr_deref_1553_Update/word_access_complete/word_0/cr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_update_start_
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1318/assign_stmt_1484_to_assign_stmt_1573/type_cast_1559_Update/cr
      -- 
    phi_stmt_1471_ack_4097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1471_ack_0, ack => convTransposeA_CP_3357_elements(87)); -- 
    rr_3624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1499_inst_req_0); -- 
    cr_3629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1499_inst_req_1); -- 
    cr_3643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1513_inst_req_1); -- 
    req_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => array_obj_ref_1519_index_offset_req_1); -- 
    req_3689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => addr_of_1520_final_reg_req_1); -- 
    cr_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => ptr_deref_1524_load_0_req_1); -- 
    rr_3748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1529_inst_req_0); -- 
    cr_3753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1529_inst_req_1); -- 
    cr_3767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1543_inst_req_1); -- 
    req_3798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => array_obj_ref_1549_index_offset_req_1); -- 
    req_3813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => addr_of_1550_final_reg_req_1); -- 
    cr_3863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => ptr_deref_1553_store_0_req_1); -- 
    rr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1559_inst_req_0); -- 
    cr_3877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3357_elements(87), ack => type_cast_1559_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1507_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1537_wire : std_logic_vector(31 downto 0);
    signal R_idxprom85_1548_resized : std_logic_vector(13 downto 0);
    signal R_idxprom85_1548_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1518_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1518_scaled : std_logic_vector(13 downto 0);
    signal add32_1489 : std_logic_vector(15 downto 0);
    signal add76_1494 : std_logic_vector(15 downto 0);
    signal add90_1566 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1519_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1519_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1519_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1519_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1519_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1519_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1549_root_address : std_logic_vector(13 downto 0);
    signal arrayidx80_1521 : std_logic_vector(31 downto 0);
    signal arrayidx86_1551 : std_logic_vector(31 downto 0);
    signal call11_1339 : std_logic_vector(15 downto 0);
    signal call13_1342 : std_logic_vector(15 downto 0);
    signal call14_1345 : std_logic_vector(15 downto 0);
    signal call15_1348 : std_logic_vector(15 downto 0);
    signal call17_1351 : std_logic_vector(15 downto 0);
    signal call19_1354 : std_logic_vector(15 downto 0);
    signal call1_1324 : std_logic_vector(15 downto 0);
    signal call3_1327 : std_logic_vector(15 downto 0);
    signal call5_1330 : std_logic_vector(15 downto 0);
    signal call7_1333 : std_logic_vector(15 downto 0);
    signal call9_1336 : std_logic_vector(15 downto 0);
    signal call_1321 : std_logic_vector(15 downto 0);
    signal cmp105_1604 : std_logic_vector(0 downto 0);
    signal cmp116_1630 : std_logic_vector(0 downto 0);
    signal cmp_1573 : std_logic_vector(0 downto 0);
    signal conv101_1599 : std_logic_vector(31 downto 0);
    signal conv104_1363 : std_logic_vector(31 downto 0);
    signal conv111_1625 : std_logic_vector(31 downto 0);
    signal conv114_1373 : std_logic_vector(31 downto 0);
    signal conv79_1500 : std_logic_vector(31 downto 0);
    signal conv83_1530 : std_logic_vector(31 downto 0);
    signal conv89_1560 : std_logic_vector(31 downto 0);
    signal conv93_1359 : std_logic_vector(31 downto 0);
    signal div115_1379 : std_logic_vector(31 downto 0);
    signal div_1369 : std_logic_vector(31 downto 0);
    signal idxprom85_1544 : std_logic_vector(63 downto 0);
    signal idxprom_1514 : std_logic_vector(63 downto 0);
    signal inc109_1608 : std_logic_vector(15 downto 0);
    signal inc109x_xinput_dim0x_x2_1613 : std_logic_vector(15 downto 0);
    signal inc_1594 : std_logic_vector(15 downto 0);
    signal indvar_1471 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1586 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1411 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1404 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1620 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1484 : std_logic_vector(15 downto 0);
    signal ptr_deref_1524_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1524_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1524_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1524_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1524_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1553_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1553_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1553_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr84_1539 : std_logic_vector(31 downto 0);
    signal shr_1509 : std_logic_vector(31 downto 0);
    signal tmp10_1468 : std_logic_vector(15 downto 0);
    signal tmp143_1423 : std_logic_vector(15 downto 0);
    signal tmp144_1428 : std_logic_vector(15 downto 0);
    signal tmp145_1433 : std_logic_vector(15 downto 0);
    signal tmp1_1390 : std_logic_vector(15 downto 0);
    signal tmp2_1438 : std_logic_vector(15 downto 0);
    signal tmp3_1443 : std_logic_vector(15 downto 0);
    signal tmp4_1396 : std_logic_vector(15 downto 0);
    signal tmp5_1401 : std_logic_vector(15 downto 0);
    signal tmp6_1448 : std_logic_vector(15 downto 0);
    signal tmp7_1453 : std_logic_vector(15 downto 0);
    signal tmp81_1525 : std_logic_vector(63 downto 0);
    signal tmp8_1458 : std_logic_vector(15 downto 0);
    signal tmp9_1463 : std_logic_vector(15 downto 0);
    signal tmp_1385 : std_logic_vector(15 downto 0);
    signal type_cast_1367_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1377_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1383_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1408_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1410_wire : std_logic_vector(15 downto 0);
    signal type_cast_1415_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1417_wire : std_logic_vector(15 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1477_wire : std_logic_vector(15 downto 0);
    signal type_cast_1482_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1498_wire : std_logic_vector(31 downto 0);
    signal type_cast_1503_wire : std_logic_vector(31 downto 0);
    signal type_cast_1506_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1512_wire : std_logic_vector(63 downto 0);
    signal type_cast_1528_wire : std_logic_vector(31 downto 0);
    signal type_cast_1533_wire : std_logic_vector(31 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1542_wire : std_logic_vector(63 downto 0);
    signal type_cast_1558_wire : std_logic_vector(31 downto 0);
    signal type_cast_1564_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1569_wire : std_logic_vector(31 downto 0);
    signal type_cast_1571_wire : std_logic_vector(31 downto 0);
    signal type_cast_1584_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1592_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1597_wire : std_logic_vector(31 downto 0);
    signal type_cast_1617_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1623_wire : std_logic_vector(31 downto 0);
    signal type_cast_1641_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1519_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1519_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1519_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1519_resized_base_address <= "00000000000000";
    array_obj_ref_1549_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1549_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1549_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1549_resized_base_address <= "00000000000000";
    ptr_deref_1524_word_offset_0 <= "00000000000000";
    ptr_deref_1553_word_offset_0 <= "00000000000000";
    type_cast_1367_wire_constant <= "00000000000000000000000000000001";
    type_cast_1377_wire_constant <= "00000000000000000000000000000001";
    type_cast_1383_wire_constant <= "1111111111111111";
    type_cast_1394_wire_constant <= "1111111111111111";
    type_cast_1408_wire_constant <= "0000000000000000";
    type_cast_1415_wire_constant <= "0000000000000000";
    type_cast_1475_wire_constant <= "0000000000000000";
    type_cast_1482_wire_constant <= "0000000000000100";
    type_cast_1506_wire_constant <= "00000000000000000000000000000010";
    type_cast_1536_wire_constant <= "00000000000000000000000000000010";
    type_cast_1564_wire_constant <= "00000000000000000000000000000100";
    type_cast_1584_wire_constant <= "0000000000000001";
    type_cast_1592_wire_constant <= "0000000000000001";
    type_cast_1617_wire_constant <= "0000000000000000";
    type_cast_1641_wire_constant <= "0000000000000001";
    phi_stmt_1404: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1408_wire_constant & type_cast_1410_wire;
      req <= phi_stmt_1404_req_0 & phi_stmt_1404_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1404",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1404_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1404,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1404
    phi_stmt_1411: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1415_wire_constant & type_cast_1417_wire;
      req <= phi_stmt_1411_req_0 & phi_stmt_1411_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1411",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1411_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1411,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1411
    phi_stmt_1471: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1475_wire_constant & type_cast_1477_wire;
      req <= phi_stmt_1471_req_0 & phi_stmt_1471_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1471",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1471_ack_0,
          idata => idata,
          odata => indvar_1471,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1471
    -- flow-through select operator MUX_1619_inst
    input_dim1x_x2_1620 <= type_cast_1617_wire_constant when (cmp105_1604(0) /=  '0') else inc_1594;
    addr_of_1520_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1520_final_reg_req_0;
      addr_of_1520_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1520_final_reg_req_1;
      addr_of_1520_final_reg_ack_1<= rack(0);
      addr_of_1520_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1520_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1519_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx80_1521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1550_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1550_final_reg_req_0;
      addr_of_1550_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1550_final_reg_req_1;
      addr_of_1550_final_reg_ack_1<= rack(0);
      addr_of_1550_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1550_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1549_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_1551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1358_inst_req_0;
      type_cast_1358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1358_inst_req_1;
      type_cast_1358_inst_ack_1<= rack(0);
      type_cast_1358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_1359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1362_inst_req_0;
      type_cast_1362_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1362_inst_req_1;
      type_cast_1362_inst_ack_1<= rack(0);
      type_cast_1362_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1362_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1363,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1372_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1372_inst_req_0;
      type_cast_1372_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1372_inst_req_1;
      type_cast_1372_inst_ack_1<= rack(0);
      type_cast_1372_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1372_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1321,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv114_1373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1410_inst_req_0;
      type_cast_1410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1410_inst_req_1;
      type_cast_1410_inst_ack_1<= rack(0);
      type_cast_1410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1410_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1417_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1417_inst_req_0;
      type_cast_1417_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1417_inst_req_1;
      type_cast_1417_inst_ack_1<= rack(0);
      type_cast_1417_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1417_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc109x_xinput_dim0x_x2_1613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1417_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1477_inst_req_0;
      type_cast_1477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1477_inst_req_1;
      type_cast_1477_inst_ack_1<= rack(0);
      type_cast_1477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1477_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1499_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1499_inst_req_0;
      type_cast_1499_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1499_inst_req_1;
      type_cast_1499_inst_ack_1<= rack(0);
      type_cast_1499_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1499_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1498_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1500,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1503_inst
    process(conv79_1500) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv79_1500(31 downto 0);
      type_cast_1503_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1508_inst
    process(ASHR_i32_i32_1507_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1507_wire(31 downto 0);
      shr_1509 <= tmp_var; -- 
    end process;
    type_cast_1513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1513_inst_req_0;
      type_cast_1513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1513_inst_req_1;
      type_cast_1513_inst_ack_1<= rack(0);
      type_cast_1513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1512_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1529_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1529_inst_req_0;
      type_cast_1529_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1529_inst_req_1;
      type_cast_1529_inst_ack_1<= rack(0);
      type_cast_1529_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1529_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1528_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1530,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1533_inst
    process(conv83_1530) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv83_1530(31 downto 0);
      type_cast_1533_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1538_inst
    process(ASHR_i32_i32_1537_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1537_wire(31 downto 0);
      shr84_1539 <= tmp_var; -- 
    end process;
    type_cast_1543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1543_inst_req_0;
      type_cast_1543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1543_inst_req_1;
      type_cast_1543_inst_ack_1<= rack(0);
      type_cast_1543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1542_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom85_1544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1559_inst_req_0;
      type_cast_1559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1559_inst_req_1;
      type_cast_1559_inst_ack_1<= rack(0);
      type_cast_1559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1558_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1569_inst
    process(add90_1566) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add90_1566(31 downto 0);
      type_cast_1569_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1571_inst
    process(conv93_1359) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv93_1359(31 downto 0);
      type_cast_1571_wire <= tmp_var; -- 
    end process;
    type_cast_1598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1598_inst_req_0;
      type_cast_1598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1598_inst_req_1;
      type_cast_1598_inst_ack_1<= rack(0);
      type_cast_1598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1597_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_1599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp105_1604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc109_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1624_inst_req_0;
      type_cast_1624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1624_inst_req_1;
      type_cast_1624_inst_ack_1<= rack(0);
      type_cast_1624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1623_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1519_index_1_rename
    process(R_idxprom_1518_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1518_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1518_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1519_index_1_resize
    process(idxprom_1514) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1514;
      ov := iv(13 downto 0);
      R_idxprom_1518_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1519_root_address_inst
    process(array_obj_ref_1519_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1519_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1519_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1549_index_1_rename
    process(R_idxprom85_1548_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom85_1548_resized;
      ov(13 downto 0) := iv;
      R_idxprom85_1548_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1549_index_1_resize
    process(idxprom85_1544) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom85_1544;
      ov := iv(13 downto 0);
      R_idxprom85_1548_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1549_root_address_inst
    process(array_obj_ref_1549_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1549_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1549_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_addr_0
    process(ptr_deref_1524_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1524_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1524_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_base_resize
    process(arrayidx80_1521) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx80_1521;
      ov := iv(13 downto 0);
      ptr_deref_1524_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_gather_scatter
    process(ptr_deref_1524_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1524_data_0;
      ov(63 downto 0) := iv;
      tmp81_1525 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1524_root_address_inst
    process(ptr_deref_1524_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1524_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1524_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_addr_0
    process(ptr_deref_1553_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1553_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1553_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_base_resize
    process(arrayidx86_1551) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx86_1551;
      ov := iv(13 downto 0);
      ptr_deref_1553_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_gather_scatter
    process(tmp81_1525) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp81_1525;
      ov(63 downto 0) := iv;
      ptr_deref_1553_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1553_root_address_inst
    process(ptr_deref_1553_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1553_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1553_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1574_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1573;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1574_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1574_branch_req_0,
          ack0 => if_stmt_1574_branch_ack_0,
          ack1 => if_stmt_1574_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1631_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp116_1630;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1631_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1631_branch_req_0,
          ack0 => if_stmt_1631_branch_ack_0,
          ack1 => if_stmt_1631_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1384_inst
    process(call9_1336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1336, type_cast_1383_wire_constant, tmp_var);
      tmp_1385 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1395_inst
    process(call7_1333) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1333, type_cast_1394_wire_constant, tmp_var);
      tmp4_1396 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1427_inst
    process(input_dim1x_x1x_xph_1404, tmp143_1423) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1404, tmp143_1423, tmp_var);
      tmp144_1428 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1442_inst
    process(tmp1_1390, tmp2_1438) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_1390, tmp2_1438, tmp_var);
      tmp3_1443 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1452_inst
    process(tmp5_1401, tmp6_1448) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1401, tmp6_1448, tmp_var);
      tmp7_1453 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1462_inst
    process(tmp3_1443, tmp8_1458) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1443, tmp8_1458, tmp_var);
      tmp9_1463 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1488_inst
    process(tmp145_1433, input_dim2x_x1_1484) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp145_1433, input_dim2x_x1_1484, tmp_var);
      add32_1489 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1493_inst
    process(tmp10_1468, input_dim2x_x1_1484) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_1468, input_dim2x_x1_1484, tmp_var);
      add76_1494 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1585_inst
    process(indvar_1471) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1471, type_cast_1584_wire_constant, tmp_var);
      indvarx_xnext_1586 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1593_inst
    process(input_dim1x_x1x_xph_1404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1404, type_cast_1592_wire_constant, tmp_var);
      inc_1594 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1612_inst
    process(inc109_1608, input_dim0x_x2x_xph_1411) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc109_1608, input_dim0x_x2x_xph_1411, tmp_var);
      inc109x_xinput_dim0x_x2_1613 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1565_inst
    process(conv89_1560) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv89_1560, type_cast_1564_wire_constant, tmp_var);
      add90_1566 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1507_inst
    process(type_cast_1503_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1503_wire, type_cast_1506_wire_constant, tmp_var);
      ASHR_i32_i32_1507_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1537_inst
    process(type_cast_1533_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1533_wire, type_cast_1536_wire_constant, tmp_var);
      ASHR_i32_i32_1537_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1603_inst
    process(conv101_1599, div_1369) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv101_1599, div_1369, tmp_var);
      cmp105_1604 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1629_inst
    process(conv111_1625, div115_1379) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv111_1625, div115_1379, tmp_var);
      cmp116_1630 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1368_inst
    process(conv104_1363) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv104_1363, type_cast_1367_wire_constant, tmp_var);
      div_1369 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1378_inst
    process(conv114_1373) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv114_1373, type_cast_1377_wire_constant, tmp_var);
      div115_1379 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1422_inst
    process(call1_1324, input_dim0x_x2x_xph_1411) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1324, input_dim0x_x2x_xph_1411, tmp_var);
      tmp143_1423 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1432_inst
    process(call3_1327, tmp144_1428) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1327, tmp144_1428, tmp_var);
      tmp145_1433 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1437_inst
    process(call13_1342, input_dim1x_x1x_xph_1404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1342, input_dim1x_x1x_xph_1404, tmp_var);
      tmp2_1438 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1447_inst
    process(call13_1342, input_dim0x_x2x_xph_1411) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1342, input_dim0x_x2x_xph_1411, tmp_var);
      tmp6_1448 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1457_inst
    process(call17_1351, tmp7_1453) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_1351, tmp7_1453, tmp_var);
      tmp8_1458 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1467_inst
    process(call19_1354, tmp9_1463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_1354, tmp9_1463, tmp_var);
      tmp10_1468 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1483_inst
    process(indvar_1471) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1471, type_cast_1482_wire_constant, tmp_var);
      input_dim2x_x1_1484 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1572_inst
    process(type_cast_1569_wire, type_cast_1571_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1569_wire, type_cast_1571_wire, tmp_var);
      cmp_1573 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1389_inst
    process(tmp_1385, call14_1345) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1385, call14_1345, tmp_var);
      tmp1_1390 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1400_inst
    process(tmp4_1396, call14_1345) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_1396, call14_1345, tmp_var);
      tmp5_1401 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1519_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1518_scaled;
      array_obj_ref_1519_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1519_index_offset_req_0;
      array_obj_ref_1519_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1519_index_offset_req_1;
      array_obj_ref_1519_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1549_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom85_1548_scaled;
      array_obj_ref_1549_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1549_index_offset_req_0;
      array_obj_ref_1549_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1549_index_offset_req_1;
      array_obj_ref_1549_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1498_inst
    process(add32_1489) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add32_1489, tmp_var);
      type_cast_1498_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1512_inst
    process(shr_1509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1509, tmp_var);
      type_cast_1512_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1528_inst
    process(add76_1494) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add76_1494, tmp_var);
      type_cast_1528_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1542_inst
    process(shr84_1539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr84_1539, tmp_var);
      type_cast_1542_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1558_inst
    process(input_dim2x_x1_1484) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1484, tmp_var);
      type_cast_1558_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1597_inst
    process(inc_1594) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1594, tmp_var);
      type_cast_1597_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1623_inst
    process(inc109x_xinput_dim0x_x2_1613) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc109x_xinput_dim0x_x2_1613, tmp_var);
      type_cast_1623_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1524_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1524_load_0_req_0;
      ptr_deref_1524_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1524_load_0_req_1;
      ptr_deref_1524_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1524_word_address_0;
      ptr_deref_1524_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1553_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1553_store_0_req_0;
      ptr_deref_1553_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1553_store_0_req_1;
      ptr_deref_1553_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1553_word_address_0;
      data_in <= ptr_deref_1553_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1344_inst RPIPE_Block0_start_1341_inst RPIPE_Block0_start_1338_inst RPIPE_Block0_start_1335_inst RPIPE_Block0_start_1347_inst RPIPE_Block0_start_1332_inst RPIPE_Block0_start_1350_inst RPIPE_Block0_start_1329_inst RPIPE_Block0_start_1326_inst RPIPE_Block0_start_1323_inst RPIPE_Block0_start_1320_inst RPIPE_Block0_start_1353_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block0_start_1344_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1341_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1338_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1335_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1347_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1332_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1350_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1329_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1326_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1323_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1320_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1353_inst_req_0;
      RPIPE_Block0_start_1344_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1341_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1338_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1335_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1347_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1332_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1350_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1329_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1326_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1323_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1320_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1353_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block0_start_1344_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1341_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1338_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1335_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1347_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1332_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1350_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1329_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1326_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1323_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1320_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1353_inst_req_1;
      RPIPE_Block0_start_1344_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1341_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1338_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1335_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1347_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1332_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1350_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1329_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1326_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1323_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1320_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1353_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call14_1345 <= data_out(191 downto 176);
      call13_1342 <= data_out(175 downto 160);
      call11_1339 <= data_out(159 downto 144);
      call9_1336 <= data_out(143 downto 128);
      call15_1348 <= data_out(127 downto 112);
      call7_1333 <= data_out(111 downto 96);
      call17_1351 <= data_out(95 downto 80);
      call5_1330 <= data_out(79 downto 64);
      call3_1327 <= data_out(63 downto 48);
      call1_1324 <= data_out(47 downto 32);
      call_1321 <= data_out(31 downto 16);
      call19_1354 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1639_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1639_inst_req_0;
      WPIPE_Block0_done_1639_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1639_inst_req_1;
      WPIPE_Block0_done_1639_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1641_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4138_start: Boolean;
  signal convTransposeB_CP_4138_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1665_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1674_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1659_inst_ack_0 : boolean;
  signal type_cast_1698_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1665_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1665_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_ack_0 : boolean;
  signal type_cast_1698_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1662_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1665_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1683_inst_req_0 : boolean;
  signal type_cast_1698_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1677_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1656_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1671_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1659_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1653_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1674_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1674_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1662_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1650_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1656_inst_ack_0 : boolean;
  signal type_cast_1702_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1662_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1662_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1677_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1683_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1683_inst_ack_1 : boolean;
  signal type_cast_1698_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1656_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1656_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1659_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_req_0 : boolean;
  signal array_obj_ref_1847_index_offset_req_0 : boolean;
  signal type_cast_1702_inst_ack_1 : boolean;
  signal type_cast_1694_inst_ack_1 : boolean;
  signal type_cast_1694_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1674_inst_req_0 : boolean;
  signal type_cast_1841_inst_req_0 : boolean;
  signal type_cast_1841_inst_ack_0 : boolean;
  signal type_cast_1827_inst_ack_0 : boolean;
  signal type_cast_1827_inst_ack_1 : boolean;
  signal type_cast_1694_inst_ack_0 : boolean;
  signal type_cast_1841_inst_req_1 : boolean;
  signal type_cast_1841_inst_ack_1 : boolean;
  signal type_cast_1827_inst_req_1 : boolean;
  signal type_cast_1694_inst_req_0 : boolean;
  signal type_cast_1827_inst_req_0 : boolean;
  signal type_cast_1702_inst_req_1 : boolean;
  signal type_cast_1702_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1683_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1659_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1650_inst_req_1 : boolean;
  signal array_obj_ref_1847_index_offset_ack_0 : boolean;
  signal array_obj_ref_1847_index_offset_req_1 : boolean;
  signal array_obj_ref_1847_index_offset_ack_1 : boolean;
  signal addr_of_1848_final_reg_req_0 : boolean;
  signal addr_of_1848_final_reg_ack_0 : boolean;
  signal addr_of_1848_final_reg_req_1 : boolean;
  signal addr_of_1848_final_reg_ack_1 : boolean;
  signal ptr_deref_1852_load_0_req_0 : boolean;
  signal ptr_deref_1852_load_0_ack_0 : boolean;
  signal ptr_deref_1852_load_0_req_1 : boolean;
  signal ptr_deref_1852_load_0_ack_1 : boolean;
  signal type_cast_1857_inst_req_0 : boolean;
  signal type_cast_1857_inst_ack_0 : boolean;
  signal type_cast_1857_inst_req_1 : boolean;
  signal type_cast_1857_inst_ack_1 : boolean;
  signal type_cast_1871_inst_req_0 : boolean;
  signal type_cast_1871_inst_ack_0 : boolean;
  signal type_cast_1871_inst_req_1 : boolean;
  signal type_cast_1871_inst_ack_1 : boolean;
  signal array_obj_ref_1877_index_offset_req_0 : boolean;
  signal array_obj_ref_1877_index_offset_ack_0 : boolean;
  signal array_obj_ref_1877_index_offset_req_1 : boolean;
  signal array_obj_ref_1877_index_offset_ack_1 : boolean;
  signal addr_of_1878_final_reg_req_0 : boolean;
  signal addr_of_1878_final_reg_ack_0 : boolean;
  signal addr_of_1878_final_reg_req_1 : boolean;
  signal addr_of_1878_final_reg_ack_1 : boolean;
  signal ptr_deref_1881_store_0_req_0 : boolean;
  signal ptr_deref_1881_store_0_ack_0 : boolean;
  signal ptr_deref_1881_store_0_req_1 : boolean;
  signal ptr_deref_1881_store_0_ack_1 : boolean;
  signal type_cast_1887_inst_req_0 : boolean;
  signal type_cast_1887_inst_ack_0 : boolean;
  signal type_cast_1887_inst_req_1 : boolean;
  signal type_cast_1887_inst_ack_1 : boolean;
  signal if_stmt_1902_branch_req_0 : boolean;
  signal if_stmt_1902_branch_ack_1 : boolean;
  signal if_stmt_1902_branch_ack_0 : boolean;
  signal type_cast_1926_inst_req_0 : boolean;
  signal type_cast_1926_inst_ack_0 : boolean;
  signal type_cast_1926_inst_req_1 : boolean;
  signal type_cast_1926_inst_ack_1 : boolean;
  signal type_cast_1941_inst_req_0 : boolean;
  signal type_cast_1941_inst_ack_0 : boolean;
  signal type_cast_1941_inst_req_1 : boolean;
  signal type_cast_1941_inst_ack_1 : boolean;
  signal type_cast_1951_inst_req_0 : boolean;
  signal type_cast_1951_inst_ack_0 : boolean;
  signal type_cast_1951_inst_req_1 : boolean;
  signal type_cast_1951_inst_ack_1 : boolean;
  signal if_stmt_1958_branch_req_0 : boolean;
  signal if_stmt_1958_branch_ack_1 : boolean;
  signal if_stmt_1958_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_1966_inst_req_0 : boolean;
  signal WPIPE_Block1_done_1966_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_1966_inst_req_1 : boolean;
  signal WPIPE_Block1_done_1966_inst_ack_1 : boolean;
  signal type_cast_1737_inst_req_0 : boolean;
  signal type_cast_1737_inst_ack_0 : boolean;
  signal type_cast_1737_inst_req_1 : boolean;
  signal type_cast_1737_inst_ack_1 : boolean;
  signal phi_stmt_1734_req_0 : boolean;
  signal phi_stmt_1740_req_0 : boolean;
  signal type_cast_1739_inst_req_0 : boolean;
  signal type_cast_1739_inst_ack_0 : boolean;
  signal type_cast_1739_inst_req_1 : boolean;
  signal type_cast_1739_inst_ack_1 : boolean;
  signal phi_stmt_1734_req_1 : boolean;
  signal type_cast_1746_inst_req_0 : boolean;
  signal type_cast_1746_inst_ack_0 : boolean;
  signal type_cast_1746_inst_req_1 : boolean;
  signal type_cast_1746_inst_ack_1 : boolean;
  signal phi_stmt_1740_req_1 : boolean;
  signal phi_stmt_1734_ack_0 : boolean;
  signal phi_stmt_1740_ack_0 : boolean;
  signal type_cast_1803_inst_req_0 : boolean;
  signal type_cast_1803_inst_ack_0 : boolean;
  signal type_cast_1803_inst_req_1 : boolean;
  signal type_cast_1803_inst_ack_1 : boolean;
  signal phi_stmt_1800_req_0 : boolean;
  signal phi_stmt_1800_req_1 : boolean;
  signal phi_stmt_1800_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4138_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4138_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4138_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4138_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4138: Block -- control-path 
    signal convTransposeB_CP_4138_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4138_elements(0) <= convTransposeB_CP_4138_start;
    convTransposeB_CP_4138_symbol <= convTransposeB_CP_4138_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1648/$entry
      -- CP-element group 0: 	 branch_block_stmt_1648/branch_block_stmt_1648__entry__
      -- CP-element group 0: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684__entry__
      -- 
    rr_4186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(0), ack => RPIPE_Block1_start_1650_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Update/cr
      -- 
    ra_4187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1650_inst_ack_0, ack => convTransposeB_CP_4138_elements(1)); -- 
    cr_4191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(1), ack => RPIPE_Block1_start_1650_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1650_Update/ca
      -- 
    ca_4192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1650_inst_ack_1, ack => convTransposeB_CP_4138_elements(2)); -- 
    rr_4200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(2), ack => RPIPE_Block1_start_1653_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_sample_completed_
      -- 
    ra_4201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1653_inst_ack_0, ack => convTransposeB_CP_4138_elements(3)); -- 
    cr_4205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(3), ack => RPIPE_Block1_start_1653_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1653_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Sample/rr
      -- 
    ca_4206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1653_inst_ack_1, ack => convTransposeB_CP_4138_elements(4)); -- 
    rr_4214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(4), ack => RPIPE_Block1_start_1656_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Update/cr
      -- 
    ra_4215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1656_inst_ack_0, ack => convTransposeB_CP_4138_elements(5)); -- 
    cr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(5), ack => RPIPE_Block1_start_1656_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1656_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Sample/$entry
      -- 
    ca_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1656_inst_ack_1, ack => convTransposeB_CP_4138_elements(6)); -- 
    rr_4228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(6), ack => RPIPE_Block1_start_1659_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Update/cr
      -- 
    ra_4229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1659_inst_ack_0, ack => convTransposeB_CP_4138_elements(7)); -- 
    cr_4233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(7), ack => RPIPE_Block1_start_1659_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1659_Update/ca
      -- 
    ca_4234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1659_inst_ack_1, ack => convTransposeB_CP_4138_elements(8)); -- 
    rr_4242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(8), ack => RPIPE_Block1_start_1662_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_sample_completed_
      -- 
    ra_4243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1662_inst_ack_0, ack => convTransposeB_CP_4138_elements(9)); -- 
    cr_4247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(9), ack => RPIPE_Block1_start_1662_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1662_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Sample/$entry
      -- 
    ca_4248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1662_inst_ack_1, ack => convTransposeB_CP_4138_elements(10)); -- 
    rr_4256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(10), ack => RPIPE_Block1_start_1665_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_update_start_
      -- 
    ra_4257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1665_inst_ack_0, ack => convTransposeB_CP_4138_elements(11)); -- 
    cr_4261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(11), ack => RPIPE_Block1_start_1665_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1665_update_completed_
      -- 
    ca_4262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1665_inst_ack_1, ack => convTransposeB_CP_4138_elements(12)); -- 
    rr_4270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(12), ack => RPIPE_Block1_start_1668_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_update_start_
      -- 
    ra_4271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1668_inst_ack_0, ack => convTransposeB_CP_4138_elements(13)); -- 
    cr_4275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(13), ack => RPIPE_Block1_start_1668_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1668_update_completed_
      -- 
    ca_4276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1668_inst_ack_1, ack => convTransposeB_CP_4138_elements(14)); -- 
    rr_4284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(14), ack => RPIPE_Block1_start_1671_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Update/cr
      -- 
    ra_4285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1671_inst_ack_0, ack => convTransposeB_CP_4138_elements(15)); -- 
    cr_4289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(15), ack => RPIPE_Block1_start_1671_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1671_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Sample/rr
      -- 
    ca_4290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1671_inst_ack_1, ack => convTransposeB_CP_4138_elements(16)); -- 
    rr_4298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(16), ack => RPIPE_Block1_start_1674_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Sample/$exit
      -- 
    ra_4299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1674_inst_ack_0, ack => convTransposeB_CP_4138_elements(17)); -- 
    cr_4303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(17), ack => RPIPE_Block1_start_1674_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1674_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_sample_start_
      -- 
    ca_4304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1674_inst_ack_1, ack => convTransposeB_CP_4138_elements(18)); -- 
    rr_4312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(18), ack => RPIPE_Block1_start_1677_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Update/cr
      -- 
    ra_4313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1677_inst_ack_0, ack => convTransposeB_CP_4138_elements(19)); -- 
    cr_4317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(19), ack => RPIPE_Block1_start_1677_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1677_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Sample/$entry
      -- 
    ca_4318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1677_inst_ack_1, ack => convTransposeB_CP_4138_elements(20)); -- 
    rr_4326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(20), ack => RPIPE_Block1_start_1680_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Update/cr
      -- 
    ra_4327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1680_inst_ack_0, ack => convTransposeB_CP_4138_elements(21)); -- 
    cr_4331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(21), ack => RPIPE_Block1_start_1680_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1680_Update/ca
      -- 
    ca_4332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1680_inst_ack_1, ack => convTransposeB_CP_4138_elements(22)); -- 
    rr_4340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(22), ack => RPIPE_Block1_start_1683_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Update/cr
      -- CP-element group 23: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Sample/ra
      -- 
    ra_4341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1683_inst_ack_0, ack => convTransposeB_CP_4138_elements(23)); -- 
    cr_4345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(23), ack => RPIPE_Block1_start_1683_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/RPIPE_Block1_start_1683_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684/$exit
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1651_to_assign_stmt_1684__exit__
      -- CP-element group 24: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731__entry__
      -- 
    ca_4346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1683_inst_ack_1, ack => convTransposeB_CP_4138_elements(24)); -- 
    rr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(24), ack => type_cast_1698_inst_req_0); -- 
    cr_4376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(24), ack => type_cast_1698_inst_req_1); -- 
    rr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(24), ack => type_cast_1702_inst_req_0); -- 
    cr_4362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(24), ack => type_cast_1694_inst_req_1); -- 
    rr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(24), ack => type_cast_1694_inst_req_0); -- 
    cr_4390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(24), ack => type_cast_1702_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Sample/$exit
      -- 
    ra_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_0, ack => convTransposeB_CP_4138_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1694_Update/$exit
      -- 
    ca_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_1, ack => convTransposeB_CP_4138_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_sample_completed_
      -- 
    ra_4372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_0, ack => convTransposeB_CP_4138_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1698_Update/ca
      -- 
    ca_4377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_1, ack => convTransposeB_CP_4138_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_sample_completed_
      -- 
    ra_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1702_inst_ack_0, ack => convTransposeB_CP_4138_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/type_cast_1702_Update/$exit
      -- 
    ca_4391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1702_inst_ack_1, ack => convTransposeB_CP_4138_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731/$exit
      -- CP-element group 31: 	 branch_block_stmt_1648/assign_stmt_1691_to_assign_stmt_1731__exit__
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/$entry
      -- CP-element group 31: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/$entry
      -- 
    rr_4781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(31), ack => type_cast_1737_inst_req_0); -- 
    cr_4786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(31), ack => type_cast_1737_inst_req_1); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(26) & convTransposeB_CP_4138_elements(28) & convTransposeB_CP_4138_elements(30);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Sample/$exit
      -- 
    ra_4406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_0, ack => convTransposeB_CP_4138_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	89 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Update/$exit
      -- 
    ca_4411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_1, ack => convTransposeB_CP_4138_elements(33)); -- 
    rr_4419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(33), ack => type_cast_1841_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Sample/$exit
      -- 
    ra_4420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1841_inst_ack_0, ack => convTransposeB_CP_4138_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	89 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_index_resize_1/index_resize_ack
      -- 
    ca_4425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1841_inst_ack_1, ack => convTransposeB_CP_4138_elements(35)); -- 
    req_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(35), ack => array_obj_ref_1847_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Sample/ack
      -- 
    ack_4451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1847_index_offset_ack_0, ack => convTransposeB_CP_4138_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	89 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_request/req
      -- 
    ack_4456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1847_index_offset_ack_1, ack => convTransposeB_CP_4138_elements(37)); -- 
    req_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(37), ack => addr_of_1848_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_request/ack
      -- 
    ack_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1848_final_reg_ack_0, ack => convTransposeB_CP_4138_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	89 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/word_access_start/word_0/rr
      -- 
    ack_4471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1848_final_reg_ack_1, ack => convTransposeB_CP_4138_elements(39)); -- 
    rr_4504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(39), ack => ptr_deref_1852_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Sample/word_access_start/word_0/ra
      -- 
    ra_4505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1852_load_0_ack_0, ack => convTransposeB_CP_4138_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	89 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/ptr_deref_1852_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/ptr_deref_1852_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/ptr_deref_1852_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/ptr_deref_1852_Merge/merge_ack
      -- 
    ca_4516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1852_load_0_ack_1, ack => convTransposeB_CP_4138_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	89 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Sample/ra
      -- 
    ra_4530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_0, ack => convTransposeB_CP_4138_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	89 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Sample/rr
      -- 
    ca_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_1, ack => convTransposeB_CP_4138_elements(43)); -- 
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(43), ack => type_cast_1871_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Sample/ra
      -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1871_inst_ack_0, ack => convTransposeB_CP_4138_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	89 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Sample/req
      -- 
    ca_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1871_inst_ack_1, ack => convTransposeB_CP_4138_elements(45)); -- 
    req_4574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(45), ack => array_obj_ref_1877_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Sample/ack
      -- 
    ack_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1877_index_offset_ack_0, ack => convTransposeB_CP_4138_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	89 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_request/req
      -- 
    ack_4580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1877_index_offset_ack_1, ack => convTransposeB_CP_4138_elements(47)); -- 
    req_4589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(47), ack => addr_of_1878_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_request/ack
      -- 
    ack_4590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1878_final_reg_ack_0, ack => convTransposeB_CP_4138_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	89 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_word_addrgen/root_register_ack
      -- 
    ack_4595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1878_final_reg_ack_1, ack => convTransposeB_CP_4138_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/ptr_deref_1881_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/ptr_deref_1881_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/ptr_deref_1881_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/ptr_deref_1881_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/word_access_start/word_0/rr
      -- 
    rr_4633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(50), ack => ptr_deref_1881_store_0_req_0); -- 
    convTransposeB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(41) & convTransposeB_CP_4138_elements(49);
      gj_convTransposeB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Sample/word_access_start/word_0/ra
      -- 
    ra_4634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1881_store_0_ack_0, ack => convTransposeB_CP_4138_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	89 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/word_access_complete/word_0/ca
      -- 
    ca_4645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1881_store_0_ack_1, ack => convTransposeB_CP_4138_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	89 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Sample/ra
      -- 
    ra_4654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1887_inst_ack_0, ack => convTransposeB_CP_4138_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	89 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Update/ca
      -- 
    ca_4659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1887_inst_ack_1, ack => convTransposeB_CP_4138_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/$exit
      -- CP-element group 55: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901__exit__
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902__entry__
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1648/R_cmp_1903_place
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1648/if_stmt_1902_else_link/$entry
      -- 
    branch_req_4667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(55), ack => if_stmt_1902_branch_req_0); -- 
    convTransposeB_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(36) & convTransposeB_CP_4138_elements(46) & convTransposeB_CP_4138_elements(52) & convTransposeB_CP_4138_elements(54);
      gj_convTransposeB_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	85 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1648/merge_stmt_1908__exit__
      -- CP-element group 56: 	 branch_block_stmt_1648/assign_stmt_1914__entry__
      -- CP-element group 56: 	 branch_block_stmt_1648/assign_stmt_1914__exit__
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1648/if_stmt_1902_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1648/if_stmt_1902_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1648/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1648/assign_stmt_1914/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/assign_stmt_1914/$exit
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1648/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1648/merge_stmt_1908_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1648/merge_stmt_1908_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1648/merge_stmt_1908_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1648/merge_stmt_1908_PhiAck/dummy
      -- 
    if_choice_transition_4672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1902_branch_ack_1, ack => convTransposeB_CP_4138_elements(56)); -- 
    rr_4870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(56), ack => type_cast_1803_inst_req_0); -- 
    cr_4875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(56), ack => type_cast_1803_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1648/merge_stmt_1916__exit__
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957__entry__
      -- CP-element group 57: 	 branch_block_stmt_1648/if_stmt_1902_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1648/if_stmt_1902_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1648/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1648/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1648/merge_stmt_1916_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1648/merge_stmt_1916_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1648/merge_stmt_1916_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1648/merge_stmt_1916_PhiAck/dummy
      -- 
    else_choice_transition_4676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1902_branch_ack_0, ack => convTransposeB_CP_4138_elements(57)); -- 
    rr_4692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(57), ack => type_cast_1926_inst_req_0); -- 
    cr_4697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(57), ack => type_cast_1926_inst_req_1); -- 
    cr_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(57), ack => type_cast_1941_inst_req_1); -- 
    cr_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(57), ack => type_cast_1951_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Sample/ra
      -- 
    ra_4693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1926_inst_ack_0, ack => convTransposeB_CP_4138_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1926_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Sample/rr
      -- 
    ca_4698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1926_inst_ack_1, ack => convTransposeB_CP_4138_elements(59)); -- 
    rr_4706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(59), ack => type_cast_1941_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Sample/ra
      -- 
    ra_4707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_0, ack => convTransposeB_CP_4138_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1941_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Sample/rr
      -- 
    ca_4712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_1, ack => convTransposeB_CP_4138_elements(61)); -- 
    rr_4720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(61), ack => type_cast_1951_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Sample/ra
      -- 
    ra_4721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_0, ack => convTransposeB_CP_4138_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957__exit__
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958__entry__
      -- CP-element group 63: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/$exit
      -- CP-element group 63: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1648/assign_stmt_1922_to_assign_stmt_1957/type_cast_1951_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1648/R_cmp132_1959_place
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1648/if_stmt_1958_else_link/$entry
      -- 
    ca_4726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1951_inst_ack_1, ack => convTransposeB_CP_4138_elements(63)); -- 
    branch_req_4734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(63), ack => if_stmt_1958_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1648/assign_stmt_1969__entry__
      -- CP-element group 64: 	 branch_block_stmt_1648/merge_stmt_1964__exit__
      -- CP-element group 64: 	 branch_block_stmt_1648/if_stmt_1958_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1648/if_stmt_1958_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1648/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1648/assign_stmt_1969/$entry
      -- CP-element group 64: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1648/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1648/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1648/merge_stmt_1964_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1648/merge_stmt_1964_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1648/merge_stmt_1964_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1648/merge_stmt_1964_PhiAck/dummy
      -- 
    if_choice_transition_4739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1958_branch_ack_1, ack => convTransposeB_CP_4138_elements(64)); -- 
    req_4756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(64), ack => WPIPE_Block1_done_1966_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	77 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1648/if_stmt_1958_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1648/if_stmt_1958_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1958_branch_ack_0, ack => convTransposeB_CP_4138_elements(65)); -- 
    rr_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(65), ack => type_cast_1739_inst_req_0); -- 
    cr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(65), ack => type_cast_1739_inst_req_1); -- 
    rr_4838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(65), ack => type_cast_1746_inst_req_0); -- 
    cr_4843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(65), ack => type_cast_1746_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Update/req
      -- 
    ack_4757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_1966_inst_ack_0, ack => convTransposeB_CP_4138_elements(66)); -- 
    req_4761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(66), ack => WPIPE_Block1_done_1966_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_1648/assign_stmt_1969__exit__
      -- CP-element group 67: 	 branch_block_stmt_1648/return__
      -- CP-element group 67: 	 branch_block_stmt_1648/merge_stmt_1971__exit__
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1648/$exit
      -- CP-element group 67: 	 branch_block_stmt_1648/branch_block_stmt_1648__exit__
      -- CP-element group 67: 	 branch_block_stmt_1648/assign_stmt_1969/$exit
      -- CP-element group 67: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1648/assign_stmt_1969/WPIPE_Block1_done_1966_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1648/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1648/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1648/merge_stmt_1971_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1648/merge_stmt_1971_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1648/merge_stmt_1971_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1648/merge_stmt_1971_PhiAck/dummy
      -- 
    ack_4762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_1966_inst_ack_1, ack => convTransposeB_CP_4138_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Sample/ra
      -- 
    ra_4782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1737_inst_ack_0, ack => convTransposeB_CP_4138_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/Update/ca
      -- 
    ca_4787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1737_inst_ack_1, ack => convTransposeB_CP_4138_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$exit
      -- CP-element group 70: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/$exit
      -- CP-element group 70: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1737/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_req
      -- 
    phi_stmt_1734_req_4788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1734_req_4788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(70), ack => phi_stmt_1734_req_0); -- 
    convTransposeB_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(68) & convTransposeB_CP_4138_elements(69);
      gj_convTransposeB_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/$exit
      -- CP-element group 71: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1744_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_req
      -- 
    phi_stmt_1740_req_4796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1740_req_4796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(71), ack => phi_stmt_1740_req_0); -- 
    -- Element group convTransposeB_CP_4138_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeB_CP_4138_elements(31), ack => convTransposeB_CP_4138_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1648/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(70) & convTransposeB_CP_4138_elements(71);
      gj_convTransposeB_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Sample/ra
      -- 
    ra_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1739_inst_ack_0, ack => convTransposeB_CP_4138_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/Update/ca
      -- 
    ca_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1739_inst_ack_1, ack => convTransposeB_CP_4138_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/$exit
      -- CP-element group 75: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/$exit
      -- CP-element group 75: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_sources/type_cast_1739/SplitProtocol/$exit
      -- CP-element group 75: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1734/phi_stmt_1734_req
      -- 
    phi_stmt_1734_req_4822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1734_req_4822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(75), ack => phi_stmt_1734_req_1); -- 
    convTransposeB_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(73) & convTransposeB_CP_4138_elements(74);
      gj_convTransposeB_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Sample/ra
      -- 
    ra_4839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1746_inst_ack_0, ack => convTransposeB_CP_4138_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/Update/ca
      -- 
    ca_4844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1746_inst_ack_1, ack => convTransposeB_CP_4138_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/$exit
      -- CP-element group 78: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/$exit
      -- CP-element group 78: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_sources/type_cast_1746/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1740/phi_stmt_1740_req
      -- 
    phi_stmt_1740_req_4845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1740_req_4845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(78), ack => phi_stmt_1740_req_1); -- 
    convTransposeB_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(76) & convTransposeB_CP_4138_elements(77);
      gj_convTransposeB_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1648/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(75) & convTransposeB_CP_4138_elements(78);
      gj_convTransposeB_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1648/merge_stmt_1733_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1648/merge_stmt_1733_PhiAck/$entry
      -- 
    convTransposeB_CP_4138_elements(80) <= OrReduce(convTransposeB_CP_4138_elements(72) & convTransposeB_CP_4138_elements(79));
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1648/merge_stmt_1733_PhiAck/phi_stmt_1734_ack
      -- 
    phi_stmt_1734_ack_4850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1734_ack_0, ack => convTransposeB_CP_4138_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1648/merge_stmt_1733_PhiAck/phi_stmt_1740_ack
      -- 
    phi_stmt_1740_ack_4851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1740_ack_0, ack => convTransposeB_CP_4138_elements(82)); -- 
    -- CP-element group 83:  join  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (10) 
      -- CP-element group 83: 	 branch_block_stmt_1648/assign_stmt_1752_to_assign_stmt_1797/$entry
      -- CP-element group 83: 	 branch_block_stmt_1648/assign_stmt_1752_to_assign_stmt_1797/$exit
      -- CP-element group 83: 	 branch_block_stmt_1648/merge_stmt_1733__exit__
      -- CP-element group 83: 	 branch_block_stmt_1648/assign_stmt_1752_to_assign_stmt_1797__entry__
      -- CP-element group 83: 	 branch_block_stmt_1648/assign_stmt_1752_to_assign_stmt_1797__exit__
      -- CP-element group 83: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 83: 	 branch_block_stmt_1648/merge_stmt_1733_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1800/$entry
      -- CP-element group 83: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$entry
      -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(81) & convTransposeB_CP_4138_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Sample/ra
      -- 
    ra_4871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_0, ack => convTransposeB_CP_4138_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/Update/ca
      -- 
    ca_4876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_1, ack => convTransposeB_CP_4138_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/$exit
      -- CP-element group 86: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/$exit
      -- CP-element group 86: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1803/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1648/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_req
      -- 
    phi_stmt_1800_req_4877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1800_req_4877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(86), ack => phi_stmt_1800_req_0); -- 
    convTransposeB_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4138_elements(84) & convTransposeB_CP_4138_elements(85);
      gj_convTransposeB_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4138_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1800/$exit
      -- CP-element group 87: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_1648/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1800/phi_stmt_1800_req
      -- 
    phi_stmt_1800_req_4888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1800_req_4888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(87), ack => phi_stmt_1800_req_1); -- 
    -- Element group convTransposeB_CP_4138_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => convTransposeB_CP_4138_elements(83), ack => convTransposeB_CP_4138_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  merge  transition  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1648/merge_stmt_1799_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1648/merge_stmt_1799_PhiAck/$entry
      -- 
    convTransposeB_CP_4138_elements(88) <= OrReduce(convTransposeB_CP_4138_elements(86) & convTransposeB_CP_4138_elements(87));
    -- CP-element group 89:  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	33 
    -- CP-element group 89: 	35 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	39 
    -- CP-element group 89: 	41 
    -- CP-element group 89: 	42 
    -- CP-element group 89: 	43 
    -- CP-element group 89: 	45 
    -- CP-element group 89: 	47 
    -- CP-element group 89: 	49 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	53 
    -- CP-element group 89: 	54 
    -- CP-element group 89:  members (51) 
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1841_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1827_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1648/merge_stmt_1799__exit__
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901__entry__
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1847_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1848_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1852_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1857_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1871_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/array_obj_ref_1877_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/addr_of_1878_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/ptr_deref_1881_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1648/assign_stmt_1813_to_assign_stmt_1901/type_cast_1887_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1648/merge_stmt_1799_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_1648/merge_stmt_1799_PhiAck/phi_stmt_1800_ack
      -- 
    phi_stmt_1800_ack_4893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1800_ack_0, ack => convTransposeB_CP_4138_elements(89)); -- 
    cr_4424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1841_inst_req_1); -- 
    cr_4410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1827_inst_req_1); -- 
    rr_4405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1827_inst_req_0); -- 
    req_4455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => array_obj_ref_1847_index_offset_req_1); -- 
    req_4470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => addr_of_1848_final_reg_req_1); -- 
    cr_4515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => ptr_deref_1852_load_0_req_1); -- 
    rr_4529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1857_inst_req_0); -- 
    cr_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1857_inst_req_1); -- 
    cr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1871_inst_req_1); -- 
    req_4579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => array_obj_ref_1877_index_offset_req_1); -- 
    req_4594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => addr_of_1878_final_reg_req_1); -- 
    cr_4644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => ptr_deref_1881_store_0_req_1); -- 
    rr_4653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1887_inst_req_0); -- 
    cr_4658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4138_elements(89), ack => type_cast_1887_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1835_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1865_wire : std_logic_vector(31 downto 0);
    signal R_idxprom96_1876_resized : std_logic_vector(13 downto 0);
    signal R_idxprom96_1876_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1846_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1846_scaled : std_logic_vector(13 downto 0);
    signal add101_1894 : std_logic_vector(31 downto 0);
    signal add43_1818 : std_logic_vector(15 downto 0);
    signal add87_1823 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1847_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1847_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1847_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1847_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1847_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1847_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1877_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1877_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1877_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1877_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1877_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1877_root_address : std_logic_vector(13 downto 0);
    signal arrayidx91_1849 : std_logic_vector(31 downto 0);
    signal arrayidx97_1879 : std_logic_vector(31 downto 0);
    signal call11_1669 : std_logic_vector(15 downto 0);
    signal call13_1672 : std_logic_vector(15 downto 0);
    signal call14_1675 : std_logic_vector(15 downto 0);
    signal call15_1678 : std_logic_vector(15 downto 0);
    signal call17_1681 : std_logic_vector(15 downto 0);
    signal call19_1684 : std_logic_vector(15 downto 0);
    signal call1_1654 : std_logic_vector(15 downto 0);
    signal call3_1657 : std_logic_vector(15 downto 0);
    signal call5_1660 : std_logic_vector(15 downto 0);
    signal call7_1663 : std_logic_vector(15 downto 0);
    signal call9_1666 : std_logic_vector(15 downto 0);
    signal call_1651 : std_logic_vector(15 downto 0);
    signal cmp116_1932 : std_logic_vector(0 downto 0);
    signal cmp132_1957 : std_logic_vector(0 downto 0);
    signal cmp_1901 : std_logic_vector(0 downto 0);
    signal conv100_1888 : std_logic_vector(31 downto 0);
    signal conv104_1695 : std_logic_vector(31 downto 0);
    signal conv112_1927 : std_logic_vector(31 downto 0);
    signal conv115_1699 : std_logic_vector(31 downto 0);
    signal conv127_1952 : std_logic_vector(31 downto 0);
    signal conv130_1703 : std_logic_vector(31 downto 0);
    signal conv90_1828 : std_logic_vector(31 downto 0);
    signal conv94_1858 : std_logic_vector(31 downto 0);
    signal div131_1709 : std_logic_vector(31 downto 0);
    signal div_1691 : std_logic_vector(15 downto 0);
    signal idxprom96_1872 : std_logic_vector(63 downto 0);
    signal idxprom_1842 : std_logic_vector(63 downto 0);
    signal inc120_1942 : std_logic_vector(15 downto 0);
    signal inc_1922 : std_logic_vector(15 downto 0);
    signal indvar_1800 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1914 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_1947 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1740 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1734 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1938 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1813 : std_logic_vector(15 downto 0);
    signal ptr_deref_1852_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1852_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1852_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1852_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1852_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1881_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1881_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1881_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1881_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1881_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1881_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr95_1867 : std_logic_vector(31 downto 0);
    signal shr_1837 : std_logic_vector(31 downto 0);
    signal tmp10_1797 : std_logic_vector(15 downto 0);
    signal tmp159_1752 : std_logic_vector(15 downto 0);
    signal tmp160_1757 : std_logic_vector(15 downto 0);
    signal tmp161_1762 : std_logic_vector(15 downto 0);
    signal tmp1_1720 : std_logic_vector(15 downto 0);
    signal tmp2_1767 : std_logic_vector(15 downto 0);
    signal tmp3_1772 : std_logic_vector(15 downto 0);
    signal tmp4_1726 : std_logic_vector(15 downto 0);
    signal tmp5_1731 : std_logic_vector(15 downto 0);
    signal tmp6_1777 : std_logic_vector(15 downto 0);
    signal tmp7_1782 : std_logic_vector(15 downto 0);
    signal tmp8_1787 : std_logic_vector(15 downto 0);
    signal tmp92_1853 : std_logic_vector(63 downto 0);
    signal tmp9_1792 : std_logic_vector(15 downto 0);
    signal tmp_1715 : std_logic_vector(15 downto 0);
    signal type_cast_1689_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1707_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1713_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1724_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1737_wire : std_logic_vector(15 downto 0);
    signal type_cast_1739_wire : std_logic_vector(15 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1746_wire : std_logic_vector(15 downto 0);
    signal type_cast_1803_wire : std_logic_vector(15 downto 0);
    signal type_cast_1806_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1811_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1826_wire : std_logic_vector(31 downto 0);
    signal type_cast_1831_wire : std_logic_vector(31 downto 0);
    signal type_cast_1834_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1840_wire : std_logic_vector(63 downto 0);
    signal type_cast_1856_wire : std_logic_vector(31 downto 0);
    signal type_cast_1861_wire : std_logic_vector(31 downto 0);
    signal type_cast_1864_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1870_wire : std_logic_vector(63 downto 0);
    signal type_cast_1886_wire : std_logic_vector(31 downto 0);
    signal type_cast_1892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1897_wire : std_logic_vector(31 downto 0);
    signal type_cast_1899_wire : std_logic_vector(31 downto 0);
    signal type_cast_1912_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1925_wire : std_logic_vector(31 downto 0);
    signal type_cast_1950_wire : std_logic_vector(31 downto 0);
    signal type_cast_1968_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1847_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1847_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1847_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1847_resized_base_address <= "00000000000000";
    array_obj_ref_1877_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1877_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1877_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1877_resized_base_address <= "00000000000000";
    ptr_deref_1852_word_offset_0 <= "00000000000000";
    ptr_deref_1881_word_offset_0 <= "00000000000000";
    type_cast_1689_wire_constant <= "0000000000000001";
    type_cast_1707_wire_constant <= "00000000000000000000000000000001";
    type_cast_1713_wire_constant <= "1111111111111111";
    type_cast_1724_wire_constant <= "1111111111111111";
    type_cast_1744_wire_constant <= "0000000000000000";
    type_cast_1806_wire_constant <= "0000000000000000";
    type_cast_1811_wire_constant <= "0000000000000100";
    type_cast_1834_wire_constant <= "00000000000000000000000000000010";
    type_cast_1864_wire_constant <= "00000000000000000000000000000010";
    type_cast_1892_wire_constant <= "00000000000000000000000000000100";
    type_cast_1912_wire_constant <= "0000000000000001";
    type_cast_1920_wire_constant <= "0000000000000001";
    type_cast_1968_wire_constant <= "0000000000000001";
    phi_stmt_1734: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1737_wire & type_cast_1739_wire;
      req <= phi_stmt_1734_req_0 & phi_stmt_1734_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1734",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1734_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1734,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1734
    phi_stmt_1740: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1744_wire_constant & type_cast_1746_wire;
      req <= phi_stmt_1740_req_0 & phi_stmt_1740_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1740",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1740_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1740,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1740
    phi_stmt_1800: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1803_wire & type_cast_1806_wire_constant;
      req <= phi_stmt_1800_req_0 & phi_stmt_1800_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1800",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1800_ack_0,
          idata => idata,
          odata => indvar_1800,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1800
    -- flow-through select operator MUX_1937_inst
    input_dim1x_x2_1938 <= div_1691 when (cmp116_1932(0) /=  '0') else inc_1922;
    addr_of_1848_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1848_final_reg_req_0;
      addr_of_1848_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1848_final_reg_req_1;
      addr_of_1848_final_reg_ack_1<= rack(0);
      addr_of_1848_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1848_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1847_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx91_1849,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1878_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1878_final_reg_req_0;
      addr_of_1878_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1878_final_reg_req_1;
      addr_of_1878_final_reg_ack_1<= rack(0);
      addr_of_1878_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1878_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1877_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx97_1879,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1694_inst_req_0;
      type_cast_1694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1694_inst_req_1;
      type_cast_1694_inst_ack_1<= rack(0);
      type_cast_1694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1657,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_1695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1698_inst_req_0;
      type_cast_1698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1698_inst_req_1;
      type_cast_1698_inst_ack_1<= rack(0);
      type_cast_1698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1699,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1702_inst_req_0;
      type_cast_1702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1702_inst_req_1;
      type_cast_1702_inst_ack_1<= rack(0);
      type_cast_1702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_1703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1737_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1737_inst_req_0;
      type_cast_1737_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1737_inst_req_1;
      type_cast_1737_inst_ack_1<= rack(0);
      type_cast_1737_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1737_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1737_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1739_inst_req_0;
      type_cast_1739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1739_inst_req_1;
      type_cast_1739_inst_ack_1<= rack(0);
      type_cast_1739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1938,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1739_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1746_inst_req_0;
      type_cast_1746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1746_inst_req_1;
      type_cast_1746_inst_ack_1<= rack(0);
      type_cast_1746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1947,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1746_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1803_inst_req_0;
      type_cast_1803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1803_inst_req_1;
      type_cast_1803_inst_ack_1<= rack(0);
      type_cast_1803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1803_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1803_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1827_inst_req_0;
      type_cast_1827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1827_inst_req_1;
      type_cast_1827_inst_ack_1<= rack(0);
      type_cast_1827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1826_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1828,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1831_inst
    process(conv90_1828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv90_1828(31 downto 0);
      type_cast_1831_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1836_inst
    process(ASHR_i32_i32_1835_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1835_wire(31 downto 0);
      shr_1837 <= tmp_var; -- 
    end process;
    type_cast_1841_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1841_inst_req_0;
      type_cast_1841_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1841_inst_req_1;
      type_cast_1841_inst_ack_1<= rack(0);
      type_cast_1841_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1841_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1840_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1842,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1857_inst_req_0;
      type_cast_1857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1857_inst_req_1;
      type_cast_1857_inst_ack_1<= rack(0);
      type_cast_1857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1856_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1861_inst
    process(conv94_1858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv94_1858(31 downto 0);
      type_cast_1861_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1866_inst
    process(ASHR_i32_i32_1865_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1865_wire(31 downto 0);
      shr95_1867 <= tmp_var; -- 
    end process;
    type_cast_1871_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1871_inst_req_0;
      type_cast_1871_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1871_inst_req_1;
      type_cast_1871_inst_ack_1<= rack(0);
      type_cast_1871_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1871_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1870_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom96_1872,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1887_inst_req_0;
      type_cast_1887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1887_inst_req_1;
      type_cast_1887_inst_ack_1<= rack(0);
      type_cast_1887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1886_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_1888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1897_inst
    process(add101_1894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add101_1894(31 downto 0);
      type_cast_1897_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1899_inst
    process(conv104_1695) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv104_1695(31 downto 0);
      type_cast_1899_wire <= tmp_var; -- 
    end process;
    type_cast_1926_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1926_inst_req_0;
      type_cast_1926_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1926_inst_req_1;
      type_cast_1926_inst_ack_1<= rack(0);
      type_cast_1926_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1926_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1925_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_1927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1941_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1941_inst_req_0;
      type_cast_1941_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1941_inst_req_1;
      type_cast_1941_inst_ack_1<= rack(0);
      type_cast_1941_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1941_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp116_1932,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc120_1942,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1951_inst_req_0;
      type_cast_1951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1951_inst_req_1;
      type_cast_1951_inst_ack_1<= rack(0);
      type_cast_1951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1950_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_1952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1847_index_1_rename
    process(R_idxprom_1846_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1846_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1846_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1847_index_1_resize
    process(idxprom_1842) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1842;
      ov := iv(13 downto 0);
      R_idxprom_1846_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1847_root_address_inst
    process(array_obj_ref_1847_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1847_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1847_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1877_index_1_rename
    process(R_idxprom96_1876_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom96_1876_resized;
      ov(13 downto 0) := iv;
      R_idxprom96_1876_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1877_index_1_resize
    process(idxprom96_1872) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom96_1872;
      ov := iv(13 downto 0);
      R_idxprom96_1876_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1877_root_address_inst
    process(array_obj_ref_1877_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1877_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1877_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1852_addr_0
    process(ptr_deref_1852_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1852_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1852_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1852_base_resize
    process(arrayidx91_1849) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx91_1849;
      ov := iv(13 downto 0);
      ptr_deref_1852_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1852_gather_scatter
    process(ptr_deref_1852_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1852_data_0;
      ov(63 downto 0) := iv;
      tmp92_1853 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1852_root_address_inst
    process(ptr_deref_1852_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1852_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1852_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1881_addr_0
    process(ptr_deref_1881_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1881_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1881_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1881_base_resize
    process(arrayidx97_1879) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx97_1879;
      ov := iv(13 downto 0);
      ptr_deref_1881_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1881_gather_scatter
    process(tmp92_1853) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp92_1853;
      ov(63 downto 0) := iv;
      ptr_deref_1881_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1881_root_address_inst
    process(ptr_deref_1881_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1881_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1881_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1902_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1901;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1902_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1902_branch_req_0,
          ack0 => if_stmt_1902_branch_ack_0,
          ack1 => if_stmt_1902_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1958_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp132_1957;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1958_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1958_branch_req_0,
          ack0 => if_stmt_1958_branch_ack_0,
          ack1 => if_stmt_1958_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1714_inst
    process(call9_1666) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1666, type_cast_1713_wire_constant, tmp_var);
      tmp_1715 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1725_inst
    process(call7_1663) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1663, type_cast_1724_wire_constant, tmp_var);
      tmp4_1726 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1756_inst
    process(input_dim1x_x1x_xph_1734, tmp159_1752) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1734, tmp159_1752, tmp_var);
      tmp160_1757 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1771_inst
    process(tmp1_1720, tmp2_1767) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_1720, tmp2_1767, tmp_var);
      tmp3_1772 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1781_inst
    process(tmp5_1731, tmp6_1777) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_1731, tmp6_1777, tmp_var);
      tmp7_1782 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1791_inst
    process(tmp3_1772, tmp8_1787) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1772, tmp8_1787, tmp_var);
      tmp9_1792 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1817_inst
    process(tmp161_1762, input_dim2x_x1_1813) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp161_1762, input_dim2x_x1_1813, tmp_var);
      add43_1818 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1822_inst
    process(tmp10_1797, input_dim2x_x1_1813) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_1797, input_dim2x_x1_1813, tmp_var);
      add87_1823 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1913_inst
    process(indvar_1800) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1800, type_cast_1912_wire_constant, tmp_var);
      indvarx_xnext_1914 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1921_inst
    process(input_dim1x_x1x_xph_1734) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1734, type_cast_1920_wire_constant, tmp_var);
      inc_1922 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1946_inst
    process(inc120_1942, input_dim0x_x2x_xph_1740) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc120_1942, input_dim0x_x2x_xph_1740, tmp_var);
      input_dim0x_x0_1947 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1893_inst
    process(conv100_1888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv100_1888, type_cast_1892_wire_constant, tmp_var);
      add101_1894 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1835_inst
    process(type_cast_1831_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1831_wire, type_cast_1834_wire_constant, tmp_var);
      ASHR_i32_i32_1835_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1865_inst
    process(type_cast_1861_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1861_wire, type_cast_1864_wire_constant, tmp_var);
      ASHR_i32_i32_1865_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1931_inst
    process(conv112_1927, conv115_1699) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_1927, conv115_1699, tmp_var);
      cmp116_1932 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1956_inst
    process(conv127_1952, div131_1709) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv127_1952, div131_1709, tmp_var);
      cmp132_1957 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1690_inst
    process(call1_1654) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call1_1654, type_cast_1689_wire_constant, tmp_var);
      div_1691 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1708_inst
    process(conv130_1703) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv130_1703, type_cast_1707_wire_constant, tmp_var);
      div131_1709 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1751_inst
    process(call1_1654, input_dim0x_x2x_xph_1740) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1654, input_dim0x_x2x_xph_1740, tmp_var);
      tmp159_1752 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1761_inst
    process(call3_1657, tmp160_1757) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1657, tmp160_1757, tmp_var);
      tmp161_1762 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1766_inst
    process(call13_1672, input_dim1x_x1x_xph_1734) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1672, input_dim1x_x1x_xph_1734, tmp_var);
      tmp2_1767 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1776_inst
    process(call13_1672, input_dim0x_x2x_xph_1740) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1672, input_dim0x_x2x_xph_1740, tmp_var);
      tmp6_1777 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1786_inst
    process(call17_1681, tmp7_1782) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_1681, tmp7_1782, tmp_var);
      tmp8_1787 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1796_inst
    process(call19_1684, tmp9_1792) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_1684, tmp9_1792, tmp_var);
      tmp10_1797 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1812_inst
    process(indvar_1800) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1800, type_cast_1811_wire_constant, tmp_var);
      input_dim2x_x1_1813 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1900_inst
    process(type_cast_1897_wire, type_cast_1899_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1897_wire, type_cast_1899_wire, tmp_var);
      cmp_1901 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1719_inst
    process(tmp_1715, call14_1675) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1715, call14_1675, tmp_var);
      tmp1_1720 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1730_inst
    process(tmp4_1726, call14_1675) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_1726, call14_1675, tmp_var);
      tmp5_1731 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1847_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1846_scaled;
      array_obj_ref_1847_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1847_index_offset_req_0;
      array_obj_ref_1847_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1847_index_offset_req_1;
      array_obj_ref_1847_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1877_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom96_1876_scaled;
      array_obj_ref_1877_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1877_index_offset_req_0;
      array_obj_ref_1877_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1877_index_offset_req_1;
      array_obj_ref_1877_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1826_inst
    process(add43_1818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add43_1818, tmp_var);
      type_cast_1826_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1840_inst
    process(shr_1837) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1837, tmp_var);
      type_cast_1840_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1856_inst
    process(add87_1823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add87_1823, tmp_var);
      type_cast_1856_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1870_inst
    process(shr95_1867) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr95_1867, tmp_var);
      type_cast_1870_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1886_inst
    process(input_dim2x_x1_1813) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1813, tmp_var);
      type_cast_1886_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1925_inst
    process(inc_1922) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1922, tmp_var);
      type_cast_1925_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1950_inst
    process(input_dim0x_x0_1947) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_1947, tmp_var);
      type_cast_1950_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1852_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1852_load_0_req_0;
      ptr_deref_1852_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1852_load_0_req_1;
      ptr_deref_1852_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1852_word_address_0;
      ptr_deref_1852_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1881_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1881_store_0_req_0;
      ptr_deref_1881_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1881_store_0_req_1;
      ptr_deref_1881_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1881_word_address_0;
      data_in <= ptr_deref_1881_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1650_inst RPIPE_Block1_start_1653_inst RPIPE_Block1_start_1656_inst RPIPE_Block1_start_1659_inst RPIPE_Block1_start_1662_inst RPIPE_Block1_start_1665_inst RPIPE_Block1_start_1668_inst RPIPE_Block1_start_1671_inst RPIPE_Block1_start_1674_inst RPIPE_Block1_start_1677_inst RPIPE_Block1_start_1680_inst RPIPE_Block1_start_1683_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_1650_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1653_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1656_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1659_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1662_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1665_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1668_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1671_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1674_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1677_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1680_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1683_inst_req_0;
      RPIPE_Block1_start_1650_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1653_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1656_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1659_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1662_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1665_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1668_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1671_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1674_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1677_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1680_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1683_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_1650_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1653_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1656_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1659_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1662_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1665_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1668_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1671_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1674_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1677_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1680_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1683_inst_req_1;
      RPIPE_Block1_start_1650_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1653_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1656_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1659_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1662_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1665_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1668_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1671_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1674_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1677_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1680_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1683_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_1651 <= data_out(191 downto 176);
      call1_1654 <= data_out(175 downto 160);
      call3_1657 <= data_out(159 downto 144);
      call5_1660 <= data_out(143 downto 128);
      call7_1663 <= data_out(127 downto 112);
      call9_1666 <= data_out(111 downto 96);
      call11_1669 <= data_out(95 downto 80);
      call13_1672 <= data_out(79 downto 64);
      call14_1675 <= data_out(63 downto 48);
      call15_1678 <= data_out(47 downto 32);
      call17_1681 <= data_out(31 downto 16);
      call19_1684 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_1966_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_1966_inst_req_0;
      WPIPE_Block1_done_1966_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_1966_inst_req_1;
      WPIPE_Block1_done_1966_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1968_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_4934_start: Boolean;
  signal convTransposeC_CP_4934_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2214_inst_req_1 : boolean;
  signal array_obj_ref_2204_index_offset_ack_0 : boolean;
  signal array_obj_ref_2174_index_offset_ack_1 : boolean;
  signal type_cast_2184_inst_ack_1 : boolean;
  signal type_cast_2262_inst_ack_1 : boolean;
  signal array_obj_ref_2174_index_offset_ack_0 : boolean;
  signal RPIPE_Block1_start_1977_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1977_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1977_inst_req_1 : boolean;
  signal type_cast_2214_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1977_inst_ack_1 : boolean;
  signal type_cast_2253_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1980_inst_req_0 : boolean;
  signal array_obj_ref_2174_index_offset_req_0 : boolean;
  signal phi_stmt_2068_req_0 : boolean;
  signal type_cast_2253_inst_req_1 : boolean;
  signal array_obj_ref_2174_index_offset_req_1 : boolean;
  signal addr_of_2175_final_reg_ack_1 : boolean;
  signal type_cast_2071_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1980_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1980_inst_req_1 : boolean;
  signal array_obj_ref_2204_index_offset_req_0 : boolean;
  signal RPIPE_Block1_start_1980_inst_ack_1 : boolean;
  signal type_cast_2071_inst_req_1 : boolean;
  signal type_cast_2214_inst_ack_1 : boolean;
  signal type_cast_2073_inst_req_1 : boolean;
  signal array_obj_ref_2204_index_offset_req_1 : boolean;
  signal array_obj_ref_2204_index_offset_ack_1 : boolean;
  signal if_stmt_2286_branch_req_0 : boolean;
  signal ptr_deref_2179_load_0_req_1 : boolean;
  signal if_stmt_2286_branch_ack_1 : boolean;
  signal ptr_deref_2179_load_0_ack_1 : boolean;
  signal if_stmt_2229_branch_req_0 : boolean;
  signal type_cast_2198_inst_req_0 : boolean;
  signal phi_stmt_2061_req_0 : boolean;
  signal addr_of_2175_final_reg_req_0 : boolean;
  signal type_cast_2279_inst_req_1 : boolean;
  signal addr_of_2205_final_reg_req_0 : boolean;
  signal type_cast_2198_inst_ack_0 : boolean;
  signal addr_of_2205_final_reg_ack_0 : boolean;
  signal if_stmt_2229_branch_ack_1 : boolean;
  signal addr_of_2175_final_reg_ack_0 : boolean;
  signal type_cast_2198_inst_req_1 : boolean;
  signal addr_of_2205_final_reg_req_1 : boolean;
  signal addr_of_2205_final_reg_ack_1 : boolean;
  signal type_cast_2073_inst_req_0 : boolean;
  signal type_cast_2184_inst_req_0 : boolean;
  signal type_cast_2184_inst_ack_0 : boolean;
  signal type_cast_2198_inst_ack_1 : boolean;
  signal type_cast_2262_inst_req_0 : boolean;
  signal if_stmt_2286_branch_ack_0 : boolean;
  signal type_cast_2073_inst_ack_0 : boolean;
  signal phi_stmt_2068_ack_0 : boolean;
  signal type_cast_2262_inst_ack_0 : boolean;
  signal type_cast_2279_inst_req_0 : boolean;
  signal type_cast_2073_inst_ack_1 : boolean;
  signal phi_stmt_2061_req_1 : boolean;
  signal type_cast_2067_inst_ack_0 : boolean;
  signal addr_of_2175_final_reg_req_1 : boolean;
  signal type_cast_2279_inst_ack_0 : boolean;
  signal phi_stmt_2061_ack_0 : boolean;
  signal if_stmt_2229_branch_ack_0 : boolean;
  signal phi_stmt_2068_req_1 : boolean;
  signal type_cast_2184_inst_req_1 : boolean;
  signal type_cast_2067_inst_req_0 : boolean;
  signal type_cast_2067_inst_req_1 : boolean;
  signal type_cast_2067_inst_ack_1 : boolean;
  signal type_cast_2214_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1983_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1983_inst_ack_0 : boolean;
  signal type_cast_2262_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1983_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1983_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1986_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1986_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1986_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1986_inst_ack_1 : boolean;
  signal type_cast_2071_inst_ack_0 : boolean;
  signal type_cast_2071_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1989_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1989_inst_ack_0 : boolean;
  signal ptr_deref_2179_load_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1989_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1989_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1992_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1992_inst_ack_0 : boolean;
  signal ptr_deref_2179_load_0_req_0 : boolean;
  signal RPIPE_Block1_start_1992_inst_req_1 : boolean;
  signal ptr_deref_2208_store_0_ack_1 : boolean;
  signal RPIPE_Block1_start_1992_inst_ack_1 : boolean;
  signal type_cast_2253_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1995_inst_req_0 : boolean;
  signal ptr_deref_2208_store_0_req_1 : boolean;
  signal RPIPE_Block1_start_1995_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1995_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1995_inst_ack_1 : boolean;
  signal type_cast_2253_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1998_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1998_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1998_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1998_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2001_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2001_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2001_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2001_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2294_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2294_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2004_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2004_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2004_inst_req_1 : boolean;
  signal ptr_deref_2208_store_0_ack_0 : boolean;
  signal RPIPE_Block1_start_2004_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2294_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2294_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2007_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2007_inst_ack_0 : boolean;
  signal ptr_deref_2208_store_0_req_0 : boolean;
  signal RPIPE_Block1_start_2007_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2007_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2010_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2010_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2010_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2010_inst_ack_1 : boolean;
  signal type_cast_2021_inst_req_0 : boolean;
  signal type_cast_2021_inst_ack_0 : boolean;
  signal type_cast_2021_inst_req_1 : boolean;
  signal type_cast_2021_inst_ack_1 : boolean;
  signal type_cast_2025_inst_req_0 : boolean;
  signal type_cast_2025_inst_ack_0 : boolean;
  signal type_cast_2279_inst_ack_1 : boolean;
  signal type_cast_2025_inst_req_1 : boolean;
  signal type_cast_2025_inst_ack_1 : boolean;
  signal type_cast_2035_inst_req_0 : boolean;
  signal type_cast_2035_inst_ack_0 : boolean;
  signal type_cast_2035_inst_req_1 : boolean;
  signal type_cast_2035_inst_ack_1 : boolean;
  signal type_cast_2154_inst_req_0 : boolean;
  signal type_cast_2154_inst_ack_0 : boolean;
  signal type_cast_2154_inst_req_1 : boolean;
  signal type_cast_2154_inst_ack_1 : boolean;
  signal type_cast_2168_inst_req_0 : boolean;
  signal type_cast_2168_inst_ack_0 : boolean;
  signal type_cast_2168_inst_req_1 : boolean;
  signal type_cast_2168_inst_ack_1 : boolean;
  signal type_cast_2133_inst_req_0 : boolean;
  signal type_cast_2133_inst_ack_0 : boolean;
  signal type_cast_2133_inst_req_1 : boolean;
  signal type_cast_2133_inst_ack_1 : boolean;
  signal phi_stmt_2127_req_1 : boolean;
  signal phi_stmt_2127_req_0 : boolean;
  signal phi_stmt_2127_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_4934_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_4934_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_4934_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_4934_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_4934: Block -- control-path 
    signal convTransposeC_CP_4934_elements: BooleanArray(89 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_4934_elements(0) <= convTransposeC_CP_4934_start;
    convTransposeC_CP_4934_symbol <= convTransposeC_CP_4934_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1975/branch_block_stmt_1975__entry__
      -- CP-element group 0: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011__entry__
      -- CP-element group 0: 	 branch_block_stmt_1975/$entry
      -- 
    rr_4982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(0), ack => RPIPE_Block1_start_1977_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_sample_completed_
      -- 
    ra_4983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1977_inst_ack_0, ack => convTransposeC_CP_4934_elements(1)); -- 
    cr_4987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(1), ack => RPIPE_Block1_start_1977_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1977_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_sample_start_
      -- 
    ca_4988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1977_inst_ack_1, ack => convTransposeC_CP_4934_elements(2)); -- 
    rr_4996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(2), ack => RPIPE_Block1_start_1980_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Update/cr
      -- 
    ra_4997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1980_inst_ack_0, ack => convTransposeC_CP_4934_elements(3)); -- 
    cr_5001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(3), ack => RPIPE_Block1_start_1980_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1980_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Sample/rr
      -- 
    ca_5002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1980_inst_ack_1, ack => convTransposeC_CP_4934_elements(4)); -- 
    rr_5010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(4), ack => RPIPE_Block1_start_1983_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Update/cr
      -- 
    ra_5011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1983_inst_ack_0, ack => convTransposeC_CP_4934_elements(5)); -- 
    cr_5015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(5), ack => RPIPE_Block1_start_1983_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1983_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Sample/rr
      -- 
    ca_5016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1983_inst_ack_1, ack => convTransposeC_CP_4934_elements(6)); -- 
    rr_5024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(6), ack => RPIPE_Block1_start_1986_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Update/cr
      -- 
    ra_5025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1986_inst_ack_0, ack => convTransposeC_CP_4934_elements(7)); -- 
    cr_5029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(7), ack => RPIPE_Block1_start_1986_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1986_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Sample/rr
      -- 
    ca_5030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1986_inst_ack_1, ack => convTransposeC_CP_4934_elements(8)); -- 
    rr_5038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(8), ack => RPIPE_Block1_start_1989_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Update/cr
      -- 
    ra_5039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1989_inst_ack_0, ack => convTransposeC_CP_4934_elements(9)); -- 
    cr_5043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(9), ack => RPIPE_Block1_start_1989_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1989_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Sample/rr
      -- 
    ca_5044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1989_inst_ack_1, ack => convTransposeC_CP_4934_elements(10)); -- 
    rr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(10), ack => RPIPE_Block1_start_1992_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Update/cr
      -- 
    ra_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1992_inst_ack_0, ack => convTransposeC_CP_4934_elements(11)); -- 
    cr_5057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(11), ack => RPIPE_Block1_start_1992_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1992_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Sample/rr
      -- 
    ca_5058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1992_inst_ack_1, ack => convTransposeC_CP_4934_elements(12)); -- 
    rr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(12), ack => RPIPE_Block1_start_1995_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Update/cr
      -- 
    ra_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1995_inst_ack_0, ack => convTransposeC_CP_4934_elements(13)); -- 
    cr_5071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(13), ack => RPIPE_Block1_start_1995_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1995_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Sample/rr
      -- 
    ca_5072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1995_inst_ack_1, ack => convTransposeC_CP_4934_elements(14)); -- 
    rr_5080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(14), ack => RPIPE_Block1_start_1998_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Update/cr
      -- 
    ra_5081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1998_inst_ack_0, ack => convTransposeC_CP_4934_elements(15)); -- 
    cr_5085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(15), ack => RPIPE_Block1_start_1998_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_1998_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Sample/rr
      -- 
    ca_5086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1998_inst_ack_1, ack => convTransposeC_CP_4934_elements(16)); -- 
    rr_5094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(16), ack => RPIPE_Block1_start_2001_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Update/cr
      -- 
    ra_5095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2001_inst_ack_0, ack => convTransposeC_CP_4934_elements(17)); -- 
    cr_5099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(17), ack => RPIPE_Block1_start_2001_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2001_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Sample/rr
      -- 
    ca_5100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2001_inst_ack_1, ack => convTransposeC_CP_4934_elements(18)); -- 
    rr_5108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(18), ack => RPIPE_Block1_start_2004_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Update/cr
      -- 
    ra_5109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2004_inst_ack_0, ack => convTransposeC_CP_4934_elements(19)); -- 
    cr_5113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(19), ack => RPIPE_Block1_start_2004_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2004_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Sample/rr
      -- 
    ca_5114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2004_inst_ack_1, ack => convTransposeC_CP_4934_elements(20)); -- 
    rr_5122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(20), ack => RPIPE_Block1_start_2007_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Update/cr
      -- 
    ra_5123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2007_inst_ack_0, ack => convTransposeC_CP_4934_elements(21)); -- 
    cr_5127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(21), ack => RPIPE_Block1_start_2007_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2007_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Sample/rr
      -- 
    ca_5128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2007_inst_ack_1, ack => convTransposeC_CP_4934_elements(22)); -- 
    rr_5136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(22), ack => RPIPE_Block1_start_2010_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Update/cr
      -- 
    ra_5137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2010_inst_ack_0, ack => convTransposeC_CP_4934_elements(23)); -- 
    cr_5141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(23), ack => RPIPE_Block1_start_2010_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011__exit__
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058__entry__
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/$exit
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_1978_to_assign_stmt_2011/RPIPE_Block1_start_2010_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Update/cr
      -- 
    ca_5142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2010_inst_ack_1, ack => convTransposeC_CP_4934_elements(24)); -- 
    rr_5153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(24), ack => type_cast_2021_inst_req_0); -- 
    cr_5158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(24), ack => type_cast_2021_inst_req_1); -- 
    rr_5167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(24), ack => type_cast_2025_inst_req_0); -- 
    cr_5172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(24), ack => type_cast_2025_inst_req_1); -- 
    rr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(24), ack => type_cast_2035_inst_req_0); -- 
    cr_5186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(24), ack => type_cast_2035_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Sample/ra
      -- 
    ra_5154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2021_inst_ack_0, ack => convTransposeC_CP_4934_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2021_Update/ca
      -- 
    ca_5159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2021_inst_ack_1, ack => convTransposeC_CP_4934_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Sample/ra
      -- 
    ra_5168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_0, ack => convTransposeC_CP_4934_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2025_Update/ca
      -- 
    ca_5173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_1, ack => convTransposeC_CP_4934_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Sample/ra
      -- 
    ra_5182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2035_inst_ack_0, ack => convTransposeC_CP_4934_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/type_cast_2035_Update/ca
      -- 
    ca_5187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2035_inst_ack_1, ack => convTransposeC_CP_4934_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058__exit__
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1975/assign_stmt_2018_to_assign_stmt_2058/$exit
      -- 
    cr_5582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(31), ack => type_cast_2071_inst_req_1); -- 
    rr_5577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(31), ack => type_cast_2071_inst_req_0); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(26) & convTransposeC_CP_4934_elements(28) & convTransposeC_CP_4934_elements(30);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	89 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Sample/ra
      -- 
    ra_5202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2154_inst_ack_0, ack => convTransposeC_CP_4934_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	89 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Sample/rr
      -- 
    ca_5207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2154_inst_ack_1, ack => convTransposeC_CP_4934_elements(33)); -- 
    rr_5215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(33), ack => type_cast_2168_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Sample/ra
      -- 
    ra_5216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2168_inst_ack_0, ack => convTransposeC_CP_4934_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	89 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Sample/req
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_index_scale_1/scale_rename_ack
      -- 
    ca_5221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2168_inst_ack_1, ack => convTransposeC_CP_4934_elements(35)); -- 
    req_5246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(35), ack => array_obj_ref_2174_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_sample_complete
      -- 
    ack_5247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2174_index_offset_ack_0, ack => convTransposeC_CP_4934_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	89 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_request/req
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_offset_calculated
      -- 
    ack_5252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2174_index_offset_ack_1, ack => convTransposeC_CP_4934_elements(37)); -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(37), ack => addr_of_2175_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_request/ack
      -- CP-element group 38: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_sample_completed_
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2175_final_reg_ack_0, ack => convTransposeC_CP_4934_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	89 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/word_access_start/word_0/rr
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_update_completed_
      -- 
    ack_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2175_final_reg_ack_1, ack => convTransposeC_CP_4934_elements(39)); -- 
    rr_5300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(39), ack => ptr_deref_2179_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/word_access_start/word_0/ra
      -- CP-element group 40: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Sample/$exit
      -- 
    ra_5301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2179_load_0_ack_0, ack => convTransposeC_CP_4934_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	89 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/ptr_deref_2179_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/ptr_deref_2179_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/ptr_deref_2179_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/ptr_deref_2179_Merge/merge_ack
      -- CP-element group 41: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_update_completed_
      -- 
    ca_5312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2179_load_0_ack_1, ack => convTransposeC_CP_4934_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	89 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Sample/ra
      -- 
    ra_5326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2184_inst_ack_0, ack => convTransposeC_CP_4934_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	89 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Update/$exit
      -- 
    ca_5331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2184_inst_ack_1, ack => convTransposeC_CP_4934_elements(43)); -- 
    rr_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(43), ack => type_cast_2198_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Sample/ra
      -- 
    ra_5340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2198_inst_ack_0, ack => convTransposeC_CP_4934_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	89 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Sample/req
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_index_resized_1
      -- 
    ca_5345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2198_inst_ack_1, ack => convTransposeC_CP_4934_elements(45)); -- 
    req_5370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(45), ack => array_obj_ref_2204_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_sample_complete
      -- 
    ack_5371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2204_index_offset_ack_0, ack => convTransposeC_CP_4934_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	89 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_request/req
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_root_address_calculated
      -- 
    ack_5376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2204_index_offset_ack_1, ack => convTransposeC_CP_4934_elements(47)); -- 
    req_5385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(47), ack => addr_of_2205_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_request/ack
      -- 
    ack_5386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2205_final_reg_ack_0, ack => convTransposeC_CP_4934_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	89 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_update_completed_
      -- 
    ack_5391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2205_final_reg_ack_1, ack => convTransposeC_CP_4934_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/ptr_deref_2208_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/word_access_start/word_0/rr
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/ptr_deref_2208_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/ptr_deref_2208_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/ptr_deref_2208_Split/$exit
      -- 
    rr_5429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(50), ack => ptr_deref_2208_store_0_req_0); -- 
    convTransposeC_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(41) & convTransposeC_CP_4934_elements(49);
      gj_convTransposeC_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/word_access_start/word_0/ra
      -- CP-element group 51: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Sample/word_access_start/$exit
      -- 
    ra_5430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2208_store_0_ack_0, ack => convTransposeC_CP_4934_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	89 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/word_access_complete/word_0/ca
      -- CP-element group 52: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/$exit
      -- 
    ca_5441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2208_store_0_ack_1, ack => convTransposeC_CP_4934_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	89 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_sample_completed_
      -- 
    ra_5450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_0, ack => convTransposeC_CP_4934_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	89 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_update_completed_
      -- 
    ca_5455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_1, ack => convTransposeC_CP_4934_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228__exit__
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229__entry__
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1975/if_stmt_2229_else_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1975/R_cmp_2230_place
      -- CP-element group 55: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/$exit
      -- 
    branch_req_5463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(55), ack => if_stmt_2229_branch_req_0); -- 
    convTransposeC_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(36) & convTransposeC_CP_4934_elements(46) & convTransposeC_CP_4934_elements(52) & convTransposeC_CP_4934_elements(54);
      gj_convTransposeC_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	85 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_1975/assign_stmt_2241__entry__
      -- CP-element group 56: 	 branch_block_stmt_1975/assign_stmt_2241__exit__
      -- CP-element group 56: 	 branch_block_stmt_1975/merge_stmt_2235__exit__
      -- CP-element group 56: 	 branch_block_stmt_1975/assign_stmt_2241/$exit
      -- CP-element group 56: 	 branch_block_stmt_1975/merge_stmt_2235_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1975/if_stmt_2229_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1975/if_stmt_2229_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/assign_stmt_2241/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1975/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1975/merge_stmt_2235_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1975/merge_stmt_2235_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1975/merge_stmt_2235_PhiAck/dummy
      -- 
    if_choice_transition_5468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2229_branch_ack_1, ack => convTransposeC_CP_4934_elements(56)); -- 
    rr_5666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(56), ack => type_cast_2133_inst_req_0); -- 
    cr_5671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(56), ack => type_cast_2133_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/merge_stmt_2243__exit__
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285__entry__
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1975/merge_stmt_2243_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1975/if_stmt_2229_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/if_stmt_2229_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1975/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1975/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1975/merge_stmt_2243_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1975/merge_stmt_2243_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1975/merge_stmt_2243_PhiAck/dummy
      -- 
    else_choice_transition_5472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2229_branch_ack_0, ack => convTransposeC_CP_4934_elements(57)); -- 
    cr_5493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(57), ack => type_cast_2253_inst_req_1); -- 
    cr_5521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(57), ack => type_cast_2279_inst_req_1); -- 
    cr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(57), ack => type_cast_2262_inst_req_1); -- 
    rr_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(57), ack => type_cast_2253_inst_req_0); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_sample_completed_
      -- 
    ra_5489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_0, ack => convTransposeC_CP_4934_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2253_update_completed_
      -- 
    ca_5494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_1, ack => convTransposeC_CP_4934_elements(59)); -- 
    rr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(59), ack => type_cast_2262_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Sample/ra
      -- 
    ra_5503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_0, ack => convTransposeC_CP_4934_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2262_Update/$exit
      -- 
    ca_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_1, ack => convTransposeC_CP_4934_elements(61)); -- 
    rr_5516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(61), ack => type_cast_2279_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Sample/$exit
      -- 
    ra_5517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_0, ack => convTransposeC_CP_4934_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285__exit__
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286__entry__
      -- CP-element group 63: 	 branch_block_stmt_1975/R_cmp128_2287_place
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286_else_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/$exit
      -- CP-element group 63: 	 branch_block_stmt_1975/if_stmt_2286_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_1975/assign_stmt_2249_to_assign_stmt_2285/type_cast_2279_Update/ca
      -- 
    ca_5522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2279_inst_ack_1, ack => convTransposeC_CP_4934_elements(63)); -- 
    branch_req_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(63), ack => if_stmt_2286_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_1975/merge_stmt_2292__exit__
      -- CP-element group 64: 	 branch_block_stmt_1975/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_1975/assign_stmt_2297__entry__
      -- CP-element group 64: 	 branch_block_stmt_1975/if_stmt_2286_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1975/if_stmt_2286_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1975/merge_stmt_2292_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1975/assign_stmt_2297/$entry
      -- CP-element group 64: 	 branch_block_stmt_1975/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1975/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1975/merge_stmt_2292_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1975/merge_stmt_2292_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1975/merge_stmt_2292_PhiAck/dummy
      -- 
    if_choice_transition_5535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2286_branch_ack_1, ack => convTransposeC_CP_4934_elements(64)); -- 
    req_5552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(64), ack => WPIPE_Block2_done_2294_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	73 
    -- CP-element group 65: 	74 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	77 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1975/if_stmt_2286_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/if_stmt_2286_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/$entry
      -- 
    else_choice_transition_5539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2286_branch_ack_0, ack => convTransposeC_CP_4934_elements(65)); -- 
    cr_5616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(65), ack => type_cast_2073_inst_req_1); -- 
    rr_5611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(65), ack => type_cast_2073_inst_req_0); -- 
    rr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(65), ack => type_cast_2067_inst_req_0); -- 
    cr_5639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(65), ack => type_cast_2067_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Update/req
      -- CP-element group 66: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_sample_completed_
      -- 
    ack_5553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2294_inst_ack_0, ack => convTransposeC_CP_4934_elements(66)); -- 
    req_5557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(66), ack => WPIPE_Block2_done_2294_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_1975/$exit
      -- CP-element group 67: 	 branch_block_stmt_1975/branch_block_stmt_1975__exit__
      -- CP-element group 67: 	 branch_block_stmt_1975/merge_stmt_2299__exit__
      -- CP-element group 67: 	 branch_block_stmt_1975/assign_stmt_2297__exit__
      -- CP-element group 67: 	 branch_block_stmt_1975/return__
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_1975/merge_stmt_2299_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1975/assign_stmt_2297/WPIPE_Block2_done_2294_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1975/assign_stmt_2297/$exit
      -- CP-element group 67: 	 branch_block_stmt_1975/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_1975/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_1975/merge_stmt_2299_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_1975/merge_stmt_2299_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_1975/merge_stmt_2299_PhiAck/dummy
      -- 
    ack_5558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2294_inst_ack_1, ack => convTransposeC_CP_4934_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Sample/ra
      -- CP-element group 68: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Sample/$exit
      -- 
    ra_5578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2071_inst_ack_0, ack => convTransposeC_CP_4934_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Update/ca
      -- CP-element group 69: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/Update/$exit
      -- 
    ca_5583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2071_inst_ack_1, ack => convTransposeC_CP_4934_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_req
      -- CP-element group 70: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2071/$exit
      -- CP-element group 70: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/$exit
      -- 
    phi_stmt_2068_req_5584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2068_req_5584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(70), ack => phi_stmt_2068_req_0); -- 
    convTransposeC_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(68) & convTransposeC_CP_4934_elements(69);
      gj_convTransposeC_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/$exit
      -- CP-element group 71: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2065_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_req
      -- 
    phi_stmt_2061_req_5592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2061_req_5592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(71), ack => phi_stmt_2061_req_0); -- 
    -- Element group convTransposeC_CP_4934_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_4934_elements(31), ack => convTransposeC_CP_4934_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  transition  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1975/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(70) & convTransposeC_CP_4934_elements(71);
      gj_convTransposeC_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	65 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Sample/ra
      -- 
    ra_5612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2073_inst_ack_0, ack => convTransposeC_CP_4934_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	65 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/Update/$exit
      -- 
    ca_5617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2073_inst_ack_1, ack => convTransposeC_CP_4934_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/$exit
      -- CP-element group 75: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/$exit
      -- CP-element group 75: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_req
      -- CP-element group 75: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2068/phi_stmt_2068_sources/type_cast_2073/SplitProtocol/$exit
      -- 
    phi_stmt_2068_req_5618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2068_req_5618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(75), ack => phi_stmt_2068_req_1); -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(73) & convTransposeC_CP_4934_elements(74);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Sample/$exit
      -- 
    ra_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_0, ack => convTransposeC_CP_4934_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	65 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/Update/ca
      -- 
    ca_5640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_1, ack => convTransposeC_CP_4934_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/$exit
      -- CP-element group 78: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_sources/type_cast_2067/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/phi_stmt_2061_req
      -- CP-element group 78: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2061/$exit
      -- 
    phi_stmt_2061_req_5641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2061_req_5641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(78), ack => phi_stmt_2061_req_1); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(76) & convTransposeC_CP_4934_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1975/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(75) & convTransposeC_CP_4934_elements(78);
      gj_convTransposeC_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1975/merge_stmt_2060_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1975/merge_stmt_2060_PhiAck/$entry
      -- 
    convTransposeC_CP_4934_elements(80) <= OrReduce(convTransposeC_CP_4934_elements(72) & convTransposeC_CP_4934_elements(79));
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1975/merge_stmt_2060_PhiAck/phi_stmt_2061_ack
      -- 
    phi_stmt_2061_ack_5646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2061_ack_0, ack => convTransposeC_CP_4934_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1975/merge_stmt_2060_PhiAck/phi_stmt_2068_ack
      -- 
    phi_stmt_2068_ack_5647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2068_ack_0, ack => convTransposeC_CP_4934_elements(82)); -- 
    -- CP-element group 83:  join  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (10) 
      -- CP-element group 83: 	 branch_block_stmt_1975/merge_stmt_2060__exit__
      -- CP-element group 83: 	 branch_block_stmt_1975/assign_stmt_2079_to_assign_stmt_2124__entry__
      -- CP-element group 83: 	 branch_block_stmt_1975/assign_stmt_2079_to_assign_stmt_2124__exit__
      -- CP-element group 83: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 83: 	 branch_block_stmt_1975/merge_stmt_2060_PhiAck/$exit
      -- CP-element group 83: 	 branch_block_stmt_1975/assign_stmt_2079_to_assign_stmt_2124/$entry
      -- CP-element group 83: 	 branch_block_stmt_1975/assign_stmt_2079_to_assign_stmt_2124/$exit
      -- CP-element group 83: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2127/$entry
      -- CP-element group 83: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/$entry
      -- 
    convTransposeC_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(81) & convTransposeC_CP_4934_elements(82);
      gj_convTransposeC_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Sample/ra
      -- 
    ra_5667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_0, ack => convTransposeC_CP_4934_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	56 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/Update/ca
      -- 
    ca_5672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2133_inst_ack_1, ack => convTransposeC_CP_4934_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/$exit
      -- CP-element group 86: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/$exit
      -- CP-element group 86: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2133/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1975/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_req
      -- 
    phi_stmt_2127_req_5673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2127_req_5673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(86), ack => phi_stmt_2127_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_4934_elements(84) & convTransposeC_CP_4934_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_4934_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  output  delay-element  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 87: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2127/$exit
      -- CP-element group 87: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_sources/type_cast_2131_konst_delay_trans
      -- CP-element group 87: 	 branch_block_stmt_1975/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2127/phi_stmt_2127_req
      -- 
    phi_stmt_2127_req_5684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2127_req_5684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(87), ack => phi_stmt_2127_req_0); -- 
    -- Element group convTransposeC_CP_4934_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => convTransposeC_CP_4934_elements(83), ack => convTransposeC_CP_4934_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  merge  transition  place  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1975/merge_stmt_2126_PhiReqMerge
      -- CP-element group 88: 	 branch_block_stmt_1975/merge_stmt_2126_PhiAck/$entry
      -- 
    convTransposeC_CP_4934_elements(88) <= OrReduce(convTransposeC_CP_4934_elements(86) & convTransposeC_CP_4934_elements(87));
    -- CP-element group 89:  fork  transition  place  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	33 
    -- CP-element group 89: 	35 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	39 
    -- CP-element group 89: 	41 
    -- CP-element group 89: 	42 
    -- CP-element group 89: 	43 
    -- CP-element group 89: 	45 
    -- CP-element group 89: 	47 
    -- CP-element group 89: 	49 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	53 
    -- CP-element group 89: 	54 
    -- CP-element group 89:  members (51) 
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228__entry__
      -- CP-element group 89: 	 branch_block_stmt_1975/merge_stmt_2126__exit__
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_Update/req
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2198_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_complete/req
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2184_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2179_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2204_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2214_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/word_access_complete/word_0/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/word_access_complete/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/word_access_complete/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/ptr_deref_2208_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2205_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2154_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/type_cast_2168_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/addr_of_2175_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1975/assign_stmt_2140_to_assign_stmt_2228/array_obj_ref_2174_final_index_sum_regn_update_start
      -- CP-element group 89: 	 branch_block_stmt_1975/merge_stmt_2126_PhiAck/$exit
      -- CP-element group 89: 	 branch_block_stmt_1975/merge_stmt_2126_PhiAck/phi_stmt_2127_ack
      -- 
    phi_stmt_2127_ack_5689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2127_ack_0, ack => convTransposeC_CP_4934_elements(89)); -- 
    cr_5454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2214_inst_req_1); -- 
    req_5251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => array_obj_ref_2174_index_offset_req_1); -- 
    req_5375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => array_obj_ref_2204_index_offset_req_1); -- 
    cr_5311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => ptr_deref_2179_load_0_req_1); -- 
    cr_5344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2198_inst_req_1); -- 
    req_5390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => addr_of_2205_final_reg_req_1); -- 
    rr_5325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2184_inst_req_0); -- 
    req_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => addr_of_2175_final_reg_req_1); -- 
    cr_5330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2184_inst_req_1); -- 
    rr_5449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2214_inst_req_0); -- 
    cr_5440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => ptr_deref_2208_store_0_req_1); -- 
    rr_5201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2154_inst_req_0); -- 
    cr_5206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2154_inst_req_1); -- 
    cr_5220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_4934_elements(89), ack => type_cast_2168_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2162_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2192_wire : std_logic_vector(31 downto 0);
    signal R_idxprom97_2203_resized : std_logic_vector(13 downto 0);
    signal R_idxprom97_2203_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2173_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2173_scaled : std_logic_vector(13 downto 0);
    signal add102_2221 : std_logic_vector(31 downto 0);
    signal add44_2145 : std_logic_vector(15 downto 0);
    signal add88_2150 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2174_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2174_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2174_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2174_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2174_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2174_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2204_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2204_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2204_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2204_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2204_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2204_root_address : std_logic_vector(13 downto 0);
    signal arrayidx92_2176 : std_logic_vector(31 downto 0);
    signal arrayidx98_2206 : std_logic_vector(31 downto 0);
    signal call11_1996 : std_logic_vector(15 downto 0);
    signal call13_1999 : std_logic_vector(15 downto 0);
    signal call14_2002 : std_logic_vector(15 downto 0);
    signal call15_2005 : std_logic_vector(15 downto 0);
    signal call17_2008 : std_logic_vector(15 downto 0);
    signal call19_2011 : std_logic_vector(15 downto 0);
    signal call1_1981 : std_logic_vector(15 downto 0);
    signal call3_1984 : std_logic_vector(15 downto 0);
    signal call5_1987 : std_logic_vector(15 downto 0);
    signal call7_1990 : std_logic_vector(15 downto 0);
    signal call9_1993 : std_logic_vector(15 downto 0);
    signal call_1978 : std_logic_vector(15 downto 0);
    signal cmp118_2259 : std_logic_vector(0 downto 0);
    signal cmp128_2285 : std_logic_vector(0 downto 0);
    signal cmp_2228 : std_logic_vector(0 downto 0);
    signal conv101_2215 : std_logic_vector(31 downto 0);
    signal conv105_2022 : std_logic_vector(31 downto 0);
    signal conv113_2254 : std_logic_vector(31 downto 0);
    signal conv116_2026 : std_logic_vector(31 downto 0);
    signal conv124_2280 : std_logic_vector(31 downto 0);
    signal conv127_2036 : std_logic_vector(31 downto 0);
    signal conv91_2155 : std_logic_vector(31 downto 0);
    signal conv95_2185 : std_logic_vector(31 downto 0);
    signal div117_2032 : std_logic_vector(31 downto 0);
    signal div_2018 : std_logic_vector(15 downto 0);
    signal idxprom97_2199 : std_logic_vector(63 downto 0);
    signal idxprom_2169 : std_logic_vector(63 downto 0);
    signal inc122_2263 : std_logic_vector(15 downto 0);
    signal inc122x_xinput_dim0x_x2_2268 : std_logic_vector(15 downto 0);
    signal inc_2249 : std_logic_vector(15 downto 0);
    signal indvar_2127 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2241 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2068 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2061 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2275 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2140 : std_logic_vector(15 downto 0);
    signal ptr_deref_2179_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2179_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2179_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2179_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2179_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2208_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2208_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2208_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2208_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2208_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2208_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr96_2194 : std_logic_vector(31 downto 0);
    signal shr_2164 : std_logic_vector(31 downto 0);
    signal tmp10_2124 : std_logic_vector(15 downto 0);
    signal tmp155_2079 : std_logic_vector(15 downto 0);
    signal tmp156_2084 : std_logic_vector(15 downto 0);
    signal tmp157_2089 : std_logic_vector(15 downto 0);
    signal tmp1_2047 : std_logic_vector(15 downto 0);
    signal tmp2_2094 : std_logic_vector(15 downto 0);
    signal tmp3_2099 : std_logic_vector(15 downto 0);
    signal tmp4_2053 : std_logic_vector(15 downto 0);
    signal tmp5_2058 : std_logic_vector(15 downto 0);
    signal tmp6_2104 : std_logic_vector(15 downto 0);
    signal tmp7_2109 : std_logic_vector(15 downto 0);
    signal tmp8_2114 : std_logic_vector(15 downto 0);
    signal tmp93_2180 : std_logic_vector(63 downto 0);
    signal tmp9_2119 : std_logic_vector(15 downto 0);
    signal tmp_2042 : std_logic_vector(15 downto 0);
    signal type_cast_2016_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2030_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2040_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2051_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2065_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2067_wire : std_logic_vector(15 downto 0);
    signal type_cast_2071_wire : std_logic_vector(15 downto 0);
    signal type_cast_2073_wire : std_logic_vector(15 downto 0);
    signal type_cast_2131_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2133_wire : std_logic_vector(15 downto 0);
    signal type_cast_2138_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2153_wire : std_logic_vector(31 downto 0);
    signal type_cast_2158_wire : std_logic_vector(31 downto 0);
    signal type_cast_2161_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2167_wire : std_logic_vector(63 downto 0);
    signal type_cast_2183_wire : std_logic_vector(31 downto 0);
    signal type_cast_2188_wire : std_logic_vector(31 downto 0);
    signal type_cast_2191_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2197_wire : std_logic_vector(63 downto 0);
    signal type_cast_2213_wire : std_logic_vector(31 downto 0);
    signal type_cast_2219_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2224_wire : std_logic_vector(31 downto 0);
    signal type_cast_2226_wire : std_logic_vector(31 downto 0);
    signal type_cast_2239_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2247_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2252_wire : std_logic_vector(31 downto 0);
    signal type_cast_2272_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2278_wire : std_logic_vector(31 downto 0);
    signal type_cast_2296_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2174_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2174_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2174_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2174_resized_base_address <= "00000000000000";
    array_obj_ref_2204_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2204_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2204_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2204_resized_base_address <= "00000000000000";
    ptr_deref_2179_word_offset_0 <= "00000000000000";
    ptr_deref_2208_word_offset_0 <= "00000000000000";
    type_cast_2016_wire_constant <= "0000000000000001";
    type_cast_2030_wire_constant <= "00000000000000000000000000000001";
    type_cast_2040_wire_constant <= "1111111111111111";
    type_cast_2051_wire_constant <= "1111111111111111";
    type_cast_2065_wire_constant <= "0000000000000000";
    type_cast_2131_wire_constant <= "0000000000000000";
    type_cast_2138_wire_constant <= "0000000000000100";
    type_cast_2161_wire_constant <= "00000000000000000000000000000010";
    type_cast_2191_wire_constant <= "00000000000000000000000000000010";
    type_cast_2219_wire_constant <= "00000000000000000000000000000100";
    type_cast_2239_wire_constant <= "0000000000000001";
    type_cast_2247_wire_constant <= "0000000000000001";
    type_cast_2272_wire_constant <= "0000000000000000";
    type_cast_2296_wire_constant <= "0000000000000001";
    phi_stmt_2061: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2065_wire_constant & type_cast_2067_wire;
      req <= phi_stmt_2061_req_0 & phi_stmt_2061_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2061",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2061_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2061,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2061
    phi_stmt_2068: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2071_wire & type_cast_2073_wire;
      req <= phi_stmt_2068_req_0 & phi_stmt_2068_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2068",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2068_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2068,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2068
    phi_stmt_2127: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2131_wire_constant & type_cast_2133_wire;
      req <= phi_stmt_2127_req_0 & phi_stmt_2127_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2127",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2127_ack_0,
          idata => idata,
          odata => indvar_2127,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2127
    -- flow-through select operator MUX_2274_inst
    input_dim1x_x2_2275 <= type_cast_2272_wire_constant when (cmp118_2259(0) /=  '0') else inc_2249;
    addr_of_2175_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2175_final_reg_req_0;
      addr_of_2175_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2175_final_reg_req_1;
      addr_of_2175_final_reg_ack_1<= rack(0);
      addr_of_2175_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2175_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2174_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2176,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2205_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2205_final_reg_req_0;
      addr_of_2205_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2205_final_reg_req_1;
      addr_of_2205_final_reg_ack_1<= rack(0);
      addr_of_2205_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2205_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2204_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx98_2206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2021_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2021_inst_req_0;
      type_cast_2021_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2021_inst_req_1;
      type_cast_2021_inst_ack_1<= rack(0);
      type_cast_2021_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2021_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv105_2022,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2025_inst_req_0;
      type_cast_2025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2025_inst_req_1;
      type_cast_2025_inst_ack_1<= rack(0);
      type_cast_2025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_1981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_2026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2035_inst_req_0;
      type_cast_2035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2035_inst_req_1;
      type_cast_2035_inst_ack_1<= rack(0);
      type_cast_2035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1978,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_2036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2067_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2067_inst_req_0;
      type_cast_2067_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2067_inst_req_1;
      type_cast_2067_inst_ack_1<= rack(0);
      type_cast_2067_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2067_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2067_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2071_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2071_inst_req_0;
      type_cast_2071_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2071_inst_req_1;
      type_cast_2071_inst_ack_1<= rack(0);
      type_cast_2071_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2071_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2071_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2073_inst_req_0;
      type_cast_2073_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2073_inst_req_1;
      type_cast_2073_inst_ack_1<= rack(0);
      type_cast_2073_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2073_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc122x_xinput_dim0x_x2_2268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2073_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2133_inst_req_0;
      type_cast_2133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2133_inst_req_1;
      type_cast_2133_inst_ack_1<= rack(0);
      type_cast_2133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2133_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2133_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2154_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2154_inst_req_0;
      type_cast_2154_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2154_inst_req_1;
      type_cast_2154_inst_ack_1<= rack(0);
      type_cast_2154_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2154_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2153_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_2155,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2158_inst
    process(conv91_2155) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv91_2155(31 downto 0);
      type_cast_2158_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2163_inst
    process(ASHR_i32_i32_2162_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2162_wire(31 downto 0);
      shr_2164 <= tmp_var; -- 
    end process;
    type_cast_2168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2168_inst_req_0;
      type_cast_2168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2168_inst_req_1;
      type_cast_2168_inst_ack_1<= rack(0);
      type_cast_2168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2167_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2184_inst_req_0;
      type_cast_2184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2184_inst_req_1;
      type_cast_2184_inst_ack_1<= rack(0);
      type_cast_2184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2183_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2185,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2188_inst
    process(conv95_2185) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv95_2185(31 downto 0);
      type_cast_2188_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2193_inst
    process(ASHR_i32_i32_2192_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2192_wire(31 downto 0);
      shr96_2194 <= tmp_var; -- 
    end process;
    type_cast_2198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2198_inst_req_0;
      type_cast_2198_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2198_inst_req_1;
      type_cast_2198_inst_ack_1<= rack(0);
      type_cast_2198_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2198_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2197_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom97_2199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2214_inst_req_0;
      type_cast_2214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2214_inst_req_1;
      type_cast_2214_inst_ack_1<= rack(0);
      type_cast_2214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2213_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_2215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2224_inst
    process(add102_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add102_2221(31 downto 0);
      type_cast_2224_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2226_inst
    process(conv105_2022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv105_2022(31 downto 0);
      type_cast_2226_wire <= tmp_var; -- 
    end process;
    type_cast_2253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2253_inst_req_0;
      type_cast_2253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2253_inst_req_1;
      type_cast_2253_inst_ack_1<= rack(0);
      type_cast_2253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2252_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_2254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2262_inst_req_0;
      type_cast_2262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2262_inst_req_1;
      type_cast_2262_inst_ack_1<= rack(0);
      type_cast_2262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp118_2259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc122_2263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2279_inst_req_0;
      type_cast_2279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2279_inst_req_1;
      type_cast_2279_inst_ack_1<= rack(0);
      type_cast_2279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2278_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv124_2280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2174_index_1_rename
    process(R_idxprom_2173_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2173_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2173_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2174_index_1_resize
    process(idxprom_2169) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2169;
      ov := iv(13 downto 0);
      R_idxprom_2173_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2174_root_address_inst
    process(array_obj_ref_2174_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2174_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2174_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2204_index_1_rename
    process(R_idxprom97_2203_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom97_2203_resized;
      ov(13 downto 0) := iv;
      R_idxprom97_2203_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2204_index_1_resize
    process(idxprom97_2199) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom97_2199;
      ov := iv(13 downto 0);
      R_idxprom97_2203_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2204_root_address_inst
    process(array_obj_ref_2204_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2204_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2204_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2179_addr_0
    process(ptr_deref_2179_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2179_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2179_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2179_base_resize
    process(arrayidx92_2176) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2176;
      ov := iv(13 downto 0);
      ptr_deref_2179_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2179_gather_scatter
    process(ptr_deref_2179_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2179_data_0;
      ov(63 downto 0) := iv;
      tmp93_2180 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2179_root_address_inst
    process(ptr_deref_2179_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2179_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2179_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2208_addr_0
    process(ptr_deref_2208_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2208_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2208_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2208_base_resize
    process(arrayidx98_2206) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx98_2206;
      ov := iv(13 downto 0);
      ptr_deref_2208_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2208_gather_scatter
    process(tmp93_2180) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp93_2180;
      ov(63 downto 0) := iv;
      ptr_deref_2208_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2208_root_address_inst
    process(ptr_deref_2208_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2208_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2208_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2229_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2228;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2229_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2229_branch_req_0,
          ack0 => if_stmt_2229_branch_ack_0,
          ack1 => if_stmt_2229_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2286_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp128_2285;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2286_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2286_branch_req_0,
          ack0 => if_stmt_2286_branch_ack_0,
          ack1 => if_stmt_2286_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2041_inst
    process(call9_1993) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1993, type_cast_2040_wire_constant, tmp_var);
      tmp_2042 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2052_inst
    process(call7_1990) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1990, type_cast_2051_wire_constant, tmp_var);
      tmp4_2053 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2083_inst
    process(input_dim1x_x1x_xph_2061, tmp155_2079) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2061, tmp155_2079, tmp_var);
      tmp156_2084 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2098_inst
    process(tmp1_2047, tmp2_2094) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_2047, tmp2_2094, tmp_var);
      tmp3_2099 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2108_inst
    process(tmp5_2058, tmp6_2104) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2058, tmp6_2104, tmp_var);
      tmp7_2109 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2118_inst
    process(tmp3_2099, tmp8_2114) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2099, tmp8_2114, tmp_var);
      tmp9_2119 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2144_inst
    process(tmp157_2089, input_dim2x_x1_2140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp157_2089, input_dim2x_x1_2140, tmp_var);
      add44_2145 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2149_inst
    process(tmp10_2124, input_dim2x_x1_2140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2124, input_dim2x_x1_2140, tmp_var);
      add88_2150 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2240_inst
    process(indvar_2127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2127, type_cast_2239_wire_constant, tmp_var);
      indvarx_xnext_2241 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2248_inst
    process(input_dim1x_x1x_xph_2061) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2061, type_cast_2247_wire_constant, tmp_var);
      inc_2249 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2267_inst
    process(inc122_2263, input_dim0x_x2x_xph_2068) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc122_2263, input_dim0x_x2x_xph_2068, tmp_var);
      inc122x_xinput_dim0x_x2_2268 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2220_inst
    process(conv101_2215) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv101_2215, type_cast_2219_wire_constant, tmp_var);
      add102_2221 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2162_inst
    process(type_cast_2158_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2158_wire, type_cast_2161_wire_constant, tmp_var);
      ASHR_i32_i32_2162_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2192_inst
    process(type_cast_2188_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2188_wire, type_cast_2191_wire_constant, tmp_var);
      ASHR_i32_i32_2192_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2258_inst
    process(conv113_2254, div117_2032) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv113_2254, div117_2032, tmp_var);
      cmp118_2259 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2284_inst
    process(conv124_2280, conv127_2036) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv124_2280, conv127_2036, tmp_var);
      cmp128_2285 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2017_inst
    process(call_1978) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1978, type_cast_2016_wire_constant, tmp_var);
      div_2018 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2031_inst
    process(conv116_2026) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv116_2026, type_cast_2030_wire_constant, tmp_var);
      div117_2032 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2078_inst
    process(call1_1981, input_dim0x_x2x_xph_2068) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_1981, input_dim0x_x2x_xph_2068, tmp_var);
      tmp155_2079 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2088_inst
    process(call3_1984, tmp156_2084) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_1984, tmp156_2084, tmp_var);
      tmp157_2089 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2093_inst
    process(call13_1999, input_dim1x_x1x_xph_2061) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1999, input_dim1x_x1x_xph_2061, tmp_var);
      tmp2_2094 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2103_inst
    process(call13_1999, input_dim0x_x2x_xph_2068) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_1999, input_dim0x_x2x_xph_2068, tmp_var);
      tmp6_2104 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2113_inst
    process(call17_2008, tmp7_2109) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_2008, tmp7_2109, tmp_var);
      tmp8_2114 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2123_inst
    process(call19_2011, tmp9_2119) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_2011, tmp9_2119, tmp_var);
      tmp10_2124 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2139_inst
    process(indvar_2127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2127, type_cast_2138_wire_constant, tmp_var);
      input_dim2x_x1_2140 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2227_inst
    process(type_cast_2224_wire, type_cast_2226_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2224_wire, type_cast_2226_wire, tmp_var);
      cmp_2228 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2046_inst
    process(tmp_2042, call14_2002) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_2042, call14_2002, tmp_var);
      tmp1_2047 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2057_inst
    process(tmp4_2053, call14_2002) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2053, call14_2002, tmp_var);
      tmp5_2058 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2174_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2173_scaled;
      array_obj_ref_2174_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2174_index_offset_req_0;
      array_obj_ref_2174_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2174_index_offset_req_1;
      array_obj_ref_2174_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2204_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom97_2203_scaled;
      array_obj_ref_2204_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2204_index_offset_req_0;
      array_obj_ref_2204_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2204_index_offset_req_1;
      array_obj_ref_2204_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2153_inst
    process(add44_2145) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add44_2145, tmp_var);
      type_cast_2153_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2167_inst
    process(shr_2164) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2164, tmp_var);
      type_cast_2167_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2183_inst
    process(add88_2150) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add88_2150, tmp_var);
      type_cast_2183_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2197_inst
    process(shr96_2194) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr96_2194, tmp_var);
      type_cast_2197_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2213_inst
    process(input_dim2x_x1_2140) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2140, tmp_var);
      type_cast_2213_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2252_inst
    process(inc_2249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2249, tmp_var);
      type_cast_2252_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2278_inst
    process(inc122x_xinput_dim0x_x2_2268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc122x_xinput_dim0x_x2_2268, tmp_var);
      type_cast_2278_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2179_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2179_load_0_req_0;
      ptr_deref_2179_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2179_load_0_req_1;
      ptr_deref_2179_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2179_word_address_0;
      ptr_deref_2179_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2208_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2208_store_0_req_0;
      ptr_deref_2208_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2208_store_0_req_1;
      ptr_deref_2208_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2208_word_address_0;
      data_in <= ptr_deref_2208_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1977_inst RPIPE_Block1_start_1980_inst RPIPE_Block1_start_1983_inst RPIPE_Block1_start_1986_inst RPIPE_Block1_start_1989_inst RPIPE_Block1_start_1992_inst RPIPE_Block1_start_1995_inst RPIPE_Block1_start_1998_inst RPIPE_Block1_start_2001_inst RPIPE_Block1_start_2004_inst RPIPE_Block1_start_2007_inst RPIPE_Block1_start_2010_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_1977_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1980_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1983_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1986_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1989_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1992_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1995_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1998_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_2001_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_2004_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_2007_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_2010_inst_req_0;
      RPIPE_Block1_start_1977_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1980_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1983_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1986_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1989_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1992_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1995_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1998_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_2001_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_2004_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_2007_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_2010_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_1977_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1980_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1983_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1986_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1989_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1992_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1995_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1998_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_2001_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_2004_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_2007_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_2010_inst_req_1;
      RPIPE_Block1_start_1977_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1980_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1983_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1986_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1989_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1992_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1995_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1998_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_2001_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_2004_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_2007_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_2010_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call_1978 <= data_out(191 downto 176);
      call1_1981 <= data_out(175 downto 160);
      call3_1984 <= data_out(159 downto 144);
      call5_1987 <= data_out(143 downto 128);
      call7_1990 <= data_out(127 downto 112);
      call9_1993 <= data_out(111 downto 96);
      call11_1996 <= data_out(95 downto 80);
      call13_1999 <= data_out(79 downto 64);
      call14_2002 <= data_out(63 downto 48);
      call15_2005 <= data_out(47 downto 32);
      call17_2008 <= data_out(31 downto 16);
      call19_2011 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2294_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2294_inst_req_0;
      WPIPE_Block2_done_2294_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2294_inst_req_1;
      WPIPE_Block2_done_2294_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2296_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_5730_start: Boolean;
  signal convTransposeD_CP_5730_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_2305_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2305_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2305_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2305_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2311_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2311_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2311_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2308_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2314_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2314_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2314_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2314_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2311_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2317_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2317_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2317_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2317_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2320_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2320_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2323_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2323_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2326_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2326_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2329_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2329_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2329_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2329_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2332_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2332_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2332_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2332_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2335_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2335_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2335_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2335_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2338_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2338_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2338_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2338_inst_ack_1 : boolean;
  signal type_cast_2355_inst_req_0 : boolean;
  signal type_cast_2355_inst_ack_0 : boolean;
  signal type_cast_2355_inst_req_1 : boolean;
  signal type_cast_2355_inst_ack_1 : boolean;
  signal type_cast_2359_inst_req_0 : boolean;
  signal type_cast_2359_inst_ack_0 : boolean;
  signal type_cast_2359_inst_req_1 : boolean;
  signal type_cast_2359_inst_ack_1 : boolean;
  signal type_cast_2363_inst_req_0 : boolean;
  signal type_cast_2363_inst_ack_0 : boolean;
  signal type_cast_2363_inst_req_1 : boolean;
  signal type_cast_2363_inst_ack_1 : boolean;
  signal type_cast_2481_inst_req_0 : boolean;
  signal type_cast_2481_inst_ack_0 : boolean;
  signal type_cast_2481_inst_req_1 : boolean;
  signal type_cast_2481_inst_ack_1 : boolean;
  signal type_cast_2495_inst_req_0 : boolean;
  signal type_cast_2495_inst_ack_0 : boolean;
  signal type_cast_2495_inst_req_1 : boolean;
  signal type_cast_2495_inst_ack_1 : boolean;
  signal array_obj_ref_2501_index_offset_req_0 : boolean;
  signal array_obj_ref_2501_index_offset_ack_0 : boolean;
  signal array_obj_ref_2501_index_offset_req_1 : boolean;
  signal array_obj_ref_2501_index_offset_ack_1 : boolean;
  signal addr_of_2502_final_reg_req_0 : boolean;
  signal addr_of_2502_final_reg_ack_0 : boolean;
  signal addr_of_2502_final_reg_req_1 : boolean;
  signal addr_of_2502_final_reg_ack_1 : boolean;
  signal ptr_deref_2506_load_0_req_0 : boolean;
  signal ptr_deref_2506_load_0_ack_0 : boolean;
  signal ptr_deref_2506_load_0_req_1 : boolean;
  signal ptr_deref_2506_load_0_ack_1 : boolean;
  signal type_cast_2511_inst_req_0 : boolean;
  signal type_cast_2511_inst_ack_0 : boolean;
  signal type_cast_2511_inst_req_1 : boolean;
  signal type_cast_2511_inst_ack_1 : boolean;
  signal type_cast_2525_inst_req_0 : boolean;
  signal type_cast_2525_inst_ack_0 : boolean;
  signal type_cast_2525_inst_req_1 : boolean;
  signal type_cast_2525_inst_ack_1 : boolean;
  signal array_obj_ref_2531_index_offset_req_0 : boolean;
  signal array_obj_ref_2531_index_offset_ack_0 : boolean;
  signal array_obj_ref_2531_index_offset_req_1 : boolean;
  signal array_obj_ref_2531_index_offset_ack_1 : boolean;
  signal addr_of_2532_final_reg_req_0 : boolean;
  signal addr_of_2532_final_reg_ack_0 : boolean;
  signal addr_of_2532_final_reg_req_1 : boolean;
  signal addr_of_2532_final_reg_ack_1 : boolean;
  signal ptr_deref_2535_store_0_req_0 : boolean;
  signal ptr_deref_2535_store_0_ack_0 : boolean;
  signal ptr_deref_2535_store_0_req_1 : boolean;
  signal ptr_deref_2535_store_0_ack_1 : boolean;
  signal type_cast_2541_inst_req_0 : boolean;
  signal type_cast_2541_inst_ack_0 : boolean;
  signal type_cast_2541_inst_req_1 : boolean;
  signal type_cast_2541_inst_ack_1 : boolean;
  signal if_stmt_2556_branch_req_0 : boolean;
  signal if_stmt_2556_branch_ack_1 : boolean;
  signal if_stmt_2556_branch_ack_0 : boolean;
  signal type_cast_2580_inst_req_0 : boolean;
  signal type_cast_2580_inst_ack_0 : boolean;
  signal type_cast_2580_inst_req_1 : boolean;
  signal type_cast_2580_inst_ack_1 : boolean;
  signal type_cast_2595_inst_req_0 : boolean;
  signal type_cast_2595_inst_ack_0 : boolean;
  signal type_cast_2595_inst_req_1 : boolean;
  signal type_cast_2595_inst_ack_1 : boolean;
  signal type_cast_2605_inst_req_0 : boolean;
  signal type_cast_2605_inst_ack_0 : boolean;
  signal type_cast_2605_inst_req_1 : boolean;
  signal type_cast_2605_inst_ack_1 : boolean;
  signal if_stmt_2612_branch_req_0 : boolean;
  signal if_stmt_2612_branch_ack_1 : boolean;
  signal if_stmt_2612_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2620_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2620_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2620_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2620_inst_ack_1 : boolean;
  signal type_cast_2394_inst_req_0 : boolean;
  signal type_cast_2394_inst_ack_0 : boolean;
  signal type_cast_2394_inst_req_1 : boolean;
  signal type_cast_2394_inst_ack_1 : boolean;
  signal phi_stmt_2389_req_1 : boolean;
  signal type_cast_2400_inst_req_0 : boolean;
  signal type_cast_2400_inst_ack_0 : boolean;
  signal type_cast_2400_inst_req_1 : boolean;
  signal type_cast_2400_inst_ack_1 : boolean;
  signal phi_stmt_2395_req_1 : boolean;
  signal type_cast_2392_inst_req_0 : boolean;
  signal type_cast_2392_inst_ack_0 : boolean;
  signal type_cast_2392_inst_req_1 : boolean;
  signal type_cast_2392_inst_ack_1 : boolean;
  signal phi_stmt_2389_req_0 : boolean;
  signal type_cast_2398_inst_req_0 : boolean;
  signal type_cast_2398_inst_ack_0 : boolean;
  signal type_cast_2398_inst_req_1 : boolean;
  signal type_cast_2398_inst_ack_1 : boolean;
  signal phi_stmt_2395_req_0 : boolean;
  signal phi_stmt_2389_ack_0 : boolean;
  signal phi_stmt_2395_ack_0 : boolean;
  signal type_cast_2457_inst_req_0 : boolean;
  signal type_cast_2457_inst_ack_0 : boolean;
  signal type_cast_2457_inst_req_1 : boolean;
  signal type_cast_2457_inst_ack_1 : boolean;
  signal phi_stmt_2454_req_0 : boolean;
  signal phi_stmt_2454_req_1 : boolean;
  signal phi_stmt_2454_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_5730_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_5730_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_5730_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_5730_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_5730: Block -- control-path 
    signal convTransposeD_CP_5730_elements: BooleanArray(91 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_5730_elements(0) <= convTransposeD_CP_5730_start;
    convTransposeD_CP_5730_symbol <= convTransposeD_CP_5730_elements(67);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2303/branch_block_stmt_2303__entry__
      -- CP-element group 0: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339__entry__
      -- CP-element group 0: 	 branch_block_stmt_2303/$entry
      -- CP-element group 0: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_5778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(0), ack => RPIPE_Block1_start_2305_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_sample_completed_
      -- 
    ra_5779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2305_inst_ack_0, ack => convTransposeD_CP_5730_elements(1)); -- 
    cr_5783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(1), ack => RPIPE_Block1_start_2305_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2305_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Sample/rr
      -- 
    ca_5784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2305_inst_ack_1, ack => convTransposeD_CP_5730_elements(2)); -- 
    rr_5792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(2), ack => RPIPE_Block1_start_2308_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Sample/$exit
      -- 
    ra_5793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2308_inst_ack_0, ack => convTransposeD_CP_5730_elements(3)); -- 
    cr_5797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(3), ack => RPIPE_Block1_start_2308_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2308_Update/$exit
      -- 
    ca_5798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2308_inst_ack_1, ack => convTransposeD_CP_5730_elements(4)); -- 
    rr_5806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(4), ack => RPIPE_Block1_start_2311_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_update_start_
      -- 
    ra_5807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2311_inst_ack_0, ack => convTransposeD_CP_5730_elements(5)); -- 
    cr_5811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(5), ack => RPIPE_Block1_start_2311_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2311_Update/ca
      -- 
    ca_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2311_inst_ack_1, ack => convTransposeD_CP_5730_elements(6)); -- 
    rr_5820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(6), ack => RPIPE_Block1_start_2314_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Sample/ra
      -- 
    ra_5821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2314_inst_ack_0, ack => convTransposeD_CP_5730_elements(7)); -- 
    cr_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(7), ack => RPIPE_Block1_start_2314_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2314_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Sample/rr
      -- 
    ca_5826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2314_inst_ack_1, ack => convTransposeD_CP_5730_elements(8)); -- 
    rr_5834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(8), ack => RPIPE_Block1_start_2317_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_update_start_
      -- CP-element group 9: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Update/cr
      -- 
    ra_5835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2317_inst_ack_0, ack => convTransposeD_CP_5730_elements(9)); -- 
    cr_5839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(9), ack => RPIPE_Block1_start_2317_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2317_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Sample/rr
      -- 
    ca_5840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2317_inst_ack_1, ack => convTransposeD_CP_5730_elements(10)); -- 
    rr_5848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(10), ack => RPIPE_Block1_start_2320_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Update/cr
      -- 
    ra_5849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2320_inst_ack_0, ack => convTransposeD_CP_5730_elements(11)); -- 
    cr_5853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(11), ack => RPIPE_Block1_start_2320_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2320_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Sample/rr
      -- 
    ca_5854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2320_inst_ack_1, ack => convTransposeD_CP_5730_elements(12)); -- 
    rr_5862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(12), ack => RPIPE_Block1_start_2323_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Update/cr
      -- 
    ra_5863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2323_inst_ack_0, ack => convTransposeD_CP_5730_elements(13)); -- 
    cr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(13), ack => RPIPE_Block1_start_2323_inst_req_1); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2323_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Sample/rr
      -- 
    ca_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2323_inst_ack_1, ack => convTransposeD_CP_5730_elements(14)); -- 
    rr_5876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(14), ack => RPIPE_Block1_start_2326_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_update_start_
      -- CP-element group 15: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Update/cr
      -- 
    ra_5877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2326_inst_ack_0, ack => convTransposeD_CP_5730_elements(15)); -- 
    cr_5881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(15), ack => RPIPE_Block1_start_2326_inst_req_1); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2326_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Sample/rr
      -- 
    ca_5882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2326_inst_ack_1, ack => convTransposeD_CP_5730_elements(16)); -- 
    rr_5890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(16), ack => RPIPE_Block1_start_2329_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_update_start_
      -- CP-element group 17: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Update/cr
      -- 
    ra_5891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2329_inst_ack_0, ack => convTransposeD_CP_5730_elements(17)); -- 
    cr_5895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(17), ack => RPIPE_Block1_start_2329_inst_req_1); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2329_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Sample/rr
      -- 
    ca_5896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2329_inst_ack_1, ack => convTransposeD_CP_5730_elements(18)); -- 
    rr_5904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(18), ack => RPIPE_Block1_start_2332_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_update_start_
      -- CP-element group 19: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Update/cr
      -- 
    ra_5905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2332_inst_ack_0, ack => convTransposeD_CP_5730_elements(19)); -- 
    cr_5909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(19), ack => RPIPE_Block1_start_2332_inst_req_1); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2332_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Sample/rr
      -- 
    ca_5910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2332_inst_ack_1, ack => convTransposeD_CP_5730_elements(20)); -- 
    rr_5918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(20), ack => RPIPE_Block1_start_2335_inst_req_0); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_update_start_
      -- CP-element group 21: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Update/cr
      -- 
    ra_5919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2335_inst_ack_0, ack => convTransposeD_CP_5730_elements(21)); -- 
    cr_5923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(21), ack => RPIPE_Block1_start_2335_inst_req_1); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2335_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Sample/rr
      -- 
    ca_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2335_inst_ack_1, ack => convTransposeD_CP_5730_elements(22)); -- 
    rr_5932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(22), ack => RPIPE_Block1_start_2338_inst_req_0); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_update_start_
      -- CP-element group 23: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Update/cr
      -- 
    ra_5933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2338_inst_ack_0, ack => convTransposeD_CP_5730_elements(23)); -- 
    cr_5937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(23), ack => RPIPE_Block1_start_2338_inst_req_1); -- 
    -- CP-element group 24:  fork  transition  place  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	29 
    -- CP-element group 24: 	30 
    -- CP-element group 24:  members (25) 
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386__entry__
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339__exit__
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/$exit
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2306_to_assign_stmt_2339/RPIPE_Block1_start_2338_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Update/cr
      -- 
    ca_5938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2338_inst_ack_1, ack => convTransposeD_CP_5730_elements(24)); -- 
    rr_5949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(24), ack => type_cast_2355_inst_req_0); -- 
    cr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(24), ack => type_cast_2355_inst_req_1); -- 
    rr_5963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(24), ack => type_cast_2359_inst_req_0); -- 
    cr_5968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(24), ack => type_cast_2359_inst_req_1); -- 
    rr_5977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(24), ack => type_cast_2363_inst_req_0); -- 
    cr_5982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(24), ack => type_cast_2363_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Sample/ra
      -- 
    ra_5950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2355_inst_ack_0, ack => convTransposeD_CP_5730_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2355_Update/ca
      -- 
    ca_5955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2355_inst_ack_1, ack => convTransposeD_CP_5730_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Sample/ra
      -- 
    ra_5964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_0, ack => convTransposeD_CP_5730_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2359_Update/ca
      -- 
    ca_5969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_1, ack => convTransposeD_CP_5730_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Sample/ra
      -- 
    ra_5978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_0, ack => convTransposeD_CP_5730_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/type_cast_2363_Update/ca
      -- 
    ca_5983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2363_inst_ack_1, ack => convTransposeD_CP_5730_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	68 
    -- CP-element group 31: 	69 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31:  members (20) 
      -- CP-element group 31: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386__exit__
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2303/assign_stmt_2346_to_assign_stmt_2386/$exit
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Update/cr
      -- 
    rr_6373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(31), ack => type_cast_2394_inst_req_0); -- 
    cr_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(31), ack => type_cast_2394_inst_req_1); -- 
    rr_6396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(31), ack => type_cast_2400_inst_req_0); -- 
    cr_6401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(31), ack => type_cast_2400_inst_req_1); -- 
    convTransposeD_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(26) & convTransposeD_CP_5730_elements(28) & convTransposeD_CP_5730_elements(30);
      gj_convTransposeD_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	91 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Sample/ra
      -- 
    ra_5998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2481_inst_ack_0, ack => convTransposeD_CP_5730_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	91 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Sample/rr
      -- 
    ca_6003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2481_inst_ack_1, ack => convTransposeD_CP_5730_elements(33)); -- 
    rr_6011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(33), ack => type_cast_2495_inst_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Sample/ra
      -- 
    ra_6012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2495_inst_ack_0, ack => convTransposeD_CP_5730_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	91 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Sample/req
      -- 
    ca_6017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2495_inst_ack_1, ack => convTransposeD_CP_5730_elements(35)); -- 
    req_6042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(35), ack => array_obj_ref_2501_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	55 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Sample/ack
      -- 
    ack_6043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2501_index_offset_ack_0, ack => convTransposeD_CP_5730_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	91 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_request/req
      -- 
    ack_6048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2501_index_offset_ack_1, ack => convTransposeD_CP_5730_elements(37)); -- 
    req_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(37), ack => addr_of_2502_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_request/ack
      -- 
    ack_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2502_final_reg_ack_0, ack => convTransposeD_CP_5730_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	91 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/word_access_start/word_0/rr
      -- 
    ack_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2502_final_reg_ack_1, ack => convTransposeD_CP_5730_elements(39)); -- 
    rr_6096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(39), ack => ptr_deref_2506_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Sample/word_access_start/word_0/ra
      -- 
    ra_6097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2506_load_0_ack_0, ack => convTransposeD_CP_5730_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	91 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/ptr_deref_2506_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/ptr_deref_2506_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/ptr_deref_2506_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/ptr_deref_2506_Merge/merge_ack
      -- 
    ca_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2506_load_0_ack_1, ack => convTransposeD_CP_5730_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	91 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Sample/ra
      -- 
    ra_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2511_inst_ack_0, ack => convTransposeD_CP_5730_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	91 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Sample/rr
      -- 
    ca_6127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2511_inst_ack_1, ack => convTransposeD_CP_5730_elements(43)); -- 
    rr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(43), ack => type_cast_2525_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Sample/ra
      -- 
    ra_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2525_inst_ack_0, ack => convTransposeD_CP_5730_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	91 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (16) 
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_resized_1
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_scaled_1
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_computed_1
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_resize_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_resize_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_resize_1/index_resize_req
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_resize_1/index_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_scale_1/$entry
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_scale_1/$exit
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_scale_1/scale_rename_req
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_index_scale_1/scale_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Sample/req
      -- 
    ca_6141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2525_inst_ack_1, ack => convTransposeD_CP_5730_elements(45)); -- 
    req_6166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(45), ack => array_obj_ref_2531_index_offset_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	55 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Sample/ack
      -- 
    ack_6167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2531_index_offset_ack_0, ack => convTransposeD_CP_5730_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	91 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_request/req
      -- 
    ack_6172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2531_index_offset_ack_1, ack => convTransposeD_CP_5730_elements(47)); -- 
    req_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(47), ack => addr_of_2532_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_request/ack
      -- 
    ack_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2532_final_reg_ack_0, ack => convTransposeD_CP_5730_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	91 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_complete/ack
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_word_addrgen/root_register_ack
      -- 
    ack_6187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2532_final_reg_ack_1, ack => convTransposeD_CP_5730_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/ptr_deref_2535_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/ptr_deref_2535_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/ptr_deref_2535_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/ptr_deref_2535_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/word_access_start/word_0/rr
      -- 
    rr_6225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(50), ack => ptr_deref_2535_store_0_req_0); -- 
    convTransposeD_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(41) & convTransposeD_CP_5730_elements(49);
      gj_convTransposeD_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Sample/word_access_start/word_0/ra
      -- 
    ra_6226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2535_store_0_ack_0, ack => convTransposeD_CP_5730_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	91 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/word_access_complete/word_0/ca
      -- 
    ca_6237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2535_store_0_ack_1, ack => convTransposeD_CP_5730_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	91 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Sample/ra
      -- 
    ra_6246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2541_inst_ack_0, ack => convTransposeD_CP_5730_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	91 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Update/ca
      -- 
    ca_6251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2541_inst_ack_1, ack => convTransposeD_CP_5730_elements(54)); -- 
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	36 
    -- CP-element group 55: 	46 
    -- CP-element group 55: 	52 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556__entry__
      -- CP-element group 55: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555__exit__
      -- CP-element group 55: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/$exit
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_2303/R_cmp_2557_place
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_2303/if_stmt_2556_else_link/$entry
      -- 
    branch_req_6259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(55), ack => if_stmt_2556_branch_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(36) & convTransposeD_CP_5730_elements(46) & convTransposeD_CP_5730_elements(52) & convTransposeD_CP_5730_elements(54);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	86 
    -- CP-element group 56: 	87 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody
      -- CP-element group 56: 	 branch_block_stmt_2303/merge_stmt_2562__exit__
      -- CP-element group 56: 	 branch_block_stmt_2303/assign_stmt_2568__exit__
      -- CP-element group 56: 	 branch_block_stmt_2303/assign_stmt_2568__entry__
      -- CP-element group 56: 	 branch_block_stmt_2303/if_stmt_2556_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_2303/if_stmt_2556_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_2303/whilex_xbody_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_2303/assign_stmt_2568/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/assign_stmt_2568/$exit
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2303/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_2303/merge_stmt_2562_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_2303/merge_stmt_2562_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_2303/merge_stmt_2562_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_2303/merge_stmt_2562_PhiAck/dummy
      -- 
    if_choice_transition_6264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2556_branch_ack_1, ack => convTransposeD_CP_5730_elements(56)); -- 
    rr_6477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(56), ack => type_cast_2457_inst_req_0); -- 
    cr_6482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(56), ack => type_cast_2457_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611__entry__
      -- CP-element group 57: 	 branch_block_stmt_2303/merge_stmt_2570__exit__
      -- CP-element group 57: 	 branch_block_stmt_2303/merge_stmt_2570_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_2303/if_stmt_2556_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_2303/if_stmt_2556_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_2303/whilex_xbody_ifx_xelse
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/$entry
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2303/merge_stmt_2570_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_update_start_
      -- CP-element group 57: 	 branch_block_stmt_2303/merge_stmt_2570_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_2303/merge_stmt_2570_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_2303/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_2303/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- 
    else_choice_transition_6268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2556_branch_ack_0, ack => convTransposeD_CP_5730_elements(57)); -- 
    rr_6284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(57), ack => type_cast_2580_inst_req_0); -- 
    cr_6289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(57), ack => type_cast_2580_inst_req_1); -- 
    cr_6303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(57), ack => type_cast_2595_inst_req_1); -- 
    cr_6317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(57), ack => type_cast_2605_inst_req_1); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Sample/ra
      -- 
    ra_6285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2580_inst_ack_0, ack => convTransposeD_CP_5730_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2580_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Sample/rr
      -- 
    ca_6290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2580_inst_ack_1, ack => convTransposeD_CP_5730_elements(59)); -- 
    rr_6298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(59), ack => type_cast_2595_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Sample/ra
      -- 
    ra_6299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2595_inst_ack_0, ack => convTransposeD_CP_5730_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2595_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Sample/rr
      -- 
    ca_6304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2595_inst_ack_1, ack => convTransposeD_CP_5730_elements(61)); -- 
    rr_6312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(61), ack => type_cast_2605_inst_req_0); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Sample/ra
      -- 
    ra_6313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2605_inst_ack_0, ack => convTransposeD_CP_5730_elements(62)); -- 
    -- CP-element group 63:  branch  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (13) 
      -- CP-element group 63: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611__exit__
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612__entry__
      -- CP-element group 63: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/$exit
      -- CP-element group 63: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2303/assign_stmt_2576_to_assign_stmt_2611/type_cast_2605_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_2303/R_cmp137_2613_place
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_2303/if_stmt_2612_else_link/$entry
      -- 
    ca_6318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2605_inst_ack_1, ack => convTransposeD_CP_5730_elements(63)); -- 
    branch_req_6326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(63), ack => if_stmt_2612_branch_req_0); -- 
    -- CP-element group 64:  merge  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (15) 
      -- CP-element group 64: 	 branch_block_stmt_2303/assign_stmt_2623__entry__
      -- CP-element group 64: 	 branch_block_stmt_2303/merge_stmt_2618__exit__
      -- CP-element group 64: 	 branch_block_stmt_2303/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_2303/merge_stmt_2618_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_2303/merge_stmt_2618_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_2303/if_stmt_2612_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_2303/merge_stmt_2618_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_2303/if_stmt_2612_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_2303/merge_stmt_2618_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_2303/ifx_xelse_whilex_xend
      -- CP-element group 64: 	 branch_block_stmt_2303/assign_stmt_2623/$entry
      -- CP-element group 64: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_2303/ifx_xelse_whilex_xend_PhiReq/$exit
      -- 
    if_choice_transition_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2612_branch_ack_1, ack => convTransposeD_CP_5730_elements(64)); -- 
    req_6348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(64), ack => WPIPE_Block3_done_2620_inst_req_0); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	75 
    -- CP-element group 65: 	76 
    -- CP-element group 65: 	78 
    -- CP-element group 65: 	79 
    -- CP-element group 65:  members (20) 
      -- CP-element group 65: 	 branch_block_stmt_2303/if_stmt_2612_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2303/if_stmt_2612_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2612_branch_ack_0, ack => convTransposeD_CP_5730_elements(65)); -- 
    rr_6422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(65), ack => type_cast_2392_inst_req_0); -- 
    cr_6427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(65), ack => type_cast_2392_inst_req_1); -- 
    rr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(65), ack => type_cast_2398_inst_req_0); -- 
    cr_6450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(65), ack => type_cast_2398_inst_req_1); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Update/req
      -- 
    ack_6349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2620_inst_ack_0, ack => convTransposeD_CP_5730_elements(66)); -- 
    req_6353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(66), ack => WPIPE_Block3_done_2620_inst_req_1); -- 
    -- CP-element group 67:  transition  place  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (16) 
      -- CP-element group 67: 	 branch_block_stmt_2303/branch_block_stmt_2303__exit__
      -- CP-element group 67: 	 $exit
      -- CP-element group 67: 	 branch_block_stmt_2303/$exit
      -- CP-element group 67: 	 branch_block_stmt_2303/merge_stmt_2625__exit__
      -- CP-element group 67: 	 branch_block_stmt_2303/return__
      -- CP-element group 67: 	 branch_block_stmt_2303/assign_stmt_2623__exit__
      -- CP-element group 67: 	 branch_block_stmt_2303/merge_stmt_2625_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2303/merge_stmt_2625_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2303/merge_stmt_2625_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2303/merge_stmt_2625_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2303/return___PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2303/return___PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2303/assign_stmt_2623/$exit
      -- CP-element group 67: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2303/assign_stmt_2623/WPIPE_Block3_done_2620_Update/ack
      -- 
    ack_6354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2620_inst_ack_1, ack => convTransposeD_CP_5730_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	31 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Sample/ra
      -- 
    ra_6374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2394_inst_ack_0, ack => convTransposeD_CP_5730_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	31 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/Update/ca
      -- 
    ca_6379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2394_inst_ack_1, ack => convTransposeD_CP_5730_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$exit
      -- CP-element group 70: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/$exit
      -- CP-element group 70: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2394/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_req
      -- 
    phi_stmt_2389_req_6380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2389_req_6380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(70), ack => phi_stmt_2389_req_1); -- 
    convTransposeD_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(68) & convTransposeD_CP_5730_elements(69);
      gj_convTransposeD_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Sample/ra
      -- 
    ra_6397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2400_inst_ack_0, ack => convTransposeD_CP_5730_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/Update/ca
      -- 
    ca_6402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2400_inst_ack_1, ack => convTransposeD_CP_5730_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/$exit
      -- CP-element group 73: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/$exit
      -- CP-element group 73: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2400/SplitProtocol/$exit
      -- CP-element group 73: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_req
      -- 
    phi_stmt_2395_req_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2395_req_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(73), ack => phi_stmt_2395_req_1); -- 
    convTransposeD_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(71) & convTransposeD_CP_5730_elements(72);
      gj_convTransposeD_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	82 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_2303/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(70) & convTransposeD_CP_5730_elements(73);
      gj_convTransposeD_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	65 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Sample/ra
      -- 
    ra_6423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2392_inst_ack_0, ack => convTransposeD_CP_5730_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	65 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/Update/ca
      -- 
    ca_6428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2392_inst_ack_1, ack => convTransposeD_CP_5730_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/$exit
      -- CP-element group 77: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/$exit
      -- CP-element group 77: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_sources/type_cast_2392/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2389/phi_stmt_2389_req
      -- 
    phi_stmt_2389_req_6429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2389_req_6429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(77), ack => phi_stmt_2389_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(75) & convTransposeD_CP_5730_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	65 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Sample/ra
      -- 
    ra_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2398_inst_ack_0, ack => convTransposeD_CP_5730_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	65 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/Update/ca
      -- 
    ca_6451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2398_inst_ack_1, ack => convTransposeD_CP_5730_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/$exit
      -- CP-element group 80: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/$exit
      -- CP-element group 80: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_sources/type_cast_2398/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2395/phi_stmt_2395_req
      -- 
    phi_stmt_2395_req_6452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2395_req_6452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(80), ack => phi_stmt_2395_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(78) & convTransposeD_CP_5730_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2303/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(77) & convTransposeD_CP_5730_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  merge  fork  transition  place  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	74 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2303/merge_stmt_2388_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_2303/merge_stmt_2388_PhiAck/$entry
      -- 
    convTransposeD_CP_5730_elements(82) <= OrReduce(convTransposeD_CP_5730_elements(74) & convTransposeD_CP_5730_elements(81));
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_2303/merge_stmt_2388_PhiAck/phi_stmt_2389_ack
      -- 
    phi_stmt_2389_ack_6457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2389_ack_0, ack => convTransposeD_CP_5730_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2303/merge_stmt_2388_PhiAck/phi_stmt_2395_ack
      -- 
    phi_stmt_2395_ack_6458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2395_ack_0, ack => convTransposeD_CP_5730_elements(84)); -- 
    -- CP-element group 85:  join  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	89 
    -- CP-element group 85:  members (10) 
      -- CP-element group 85: 	 branch_block_stmt_2303/assign_stmt_2406_to_assign_stmt_2451__exit__
      -- CP-element group 85: 	 branch_block_stmt_2303/assign_stmt_2406_to_assign_stmt_2451__entry__
      -- CP-element group 85: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 85: 	 branch_block_stmt_2303/merge_stmt_2388__exit__
      -- CP-element group 85: 	 branch_block_stmt_2303/assign_stmt_2406_to_assign_stmt_2451/$entry
      -- CP-element group 85: 	 branch_block_stmt_2303/assign_stmt_2406_to_assign_stmt_2451/$exit
      -- CP-element group 85: 	 branch_block_stmt_2303/merge_stmt_2388_PhiAck/$exit
      -- CP-element group 85: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2454/$entry
      -- CP-element group 85: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/$entry
      -- 
    convTransposeD_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(83) & convTransposeD_CP_5730_elements(84);
      gj_convTransposeD_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	56 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Sample/ra
      -- 
    ra_6478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2457_inst_ack_0, ack => convTransposeD_CP_5730_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	56 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/Update/ca
      -- 
    ca_6483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2457_inst_ack_1, ack => convTransposeD_CP_5730_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 88: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/$exit
      -- CP-element group 88: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/$exit
      -- CP-element group 88: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2457/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2303/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_req
      -- 
    phi_stmt_2454_req_6484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2454_req_6484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(88), ack => phi_stmt_2454_req_0); -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_5730_elements(86) & convTransposeD_CP_5730_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_5730_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	85 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2454/$exit
      -- CP-element group 89: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_sources/type_cast_2460_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_2303/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2454/phi_stmt_2454_req
      -- 
    phi_stmt_2454_req_6495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2454_req_6495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(89), ack => phi_stmt_2454_req_1); -- 
    -- Element group convTransposeD_CP_5730_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => convTransposeD_CP_5730_elements(85), ack => convTransposeD_CP_5730_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  merge  transition  place  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2303/merge_stmt_2453_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_2303/merge_stmt_2453_PhiAck/$entry
      -- 
    convTransposeD_CP_5730_elements(90) <= OrReduce(convTransposeD_CP_5730_elements(88) & convTransposeD_CP_5730_elements(89));
    -- CP-element group 91:  fork  transition  place  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	32 
    -- CP-element group 91: 	33 
    -- CP-element group 91: 	35 
    -- CP-element group 91: 	37 
    -- CP-element group 91: 	39 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	42 
    -- CP-element group 91: 	43 
    -- CP-element group 91: 	45 
    -- CP-element group 91: 	47 
    -- CP-element group 91: 	49 
    -- CP-element group 91: 	52 
    -- CP-element group 91: 	53 
    -- CP-element group 91: 	54 
    -- CP-element group 91:  members (51) 
      -- CP-element group 91: 	 branch_block_stmt_2303/merge_stmt_2453__exit__
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555__entry__
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2481_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2495_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_update_start
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2501_final_index_sum_regn_Update/req
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2502_complete/req
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2506_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2511_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2525_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_update_start
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/array_obj_ref_2531_final_index_sum_regn_Update/req
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/addr_of_2532_complete/req
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/word_access_complete/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/word_access_complete/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/ptr_deref_2535_Update/word_access_complete/word_0/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2303/assign_stmt_2467_to_assign_stmt_2555/type_cast_2541_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_2303/merge_stmt_2453_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_2303/merge_stmt_2453_PhiAck/phi_stmt_2454_ack
      -- 
    phi_stmt_2454_ack_6500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2454_ack_0, ack => convTransposeD_CP_5730_elements(91)); -- 
    rr_5997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2481_inst_req_0); -- 
    cr_6002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2481_inst_req_1); -- 
    cr_6016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2495_inst_req_1); -- 
    req_6047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => array_obj_ref_2501_index_offset_req_1); -- 
    req_6062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => addr_of_2502_final_reg_req_1); -- 
    cr_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => ptr_deref_2506_load_0_req_1); -- 
    rr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2511_inst_req_0); -- 
    cr_6126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2511_inst_req_1); -- 
    cr_6140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2525_inst_req_1); -- 
    req_6171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => array_obj_ref_2531_index_offset_req_1); -- 
    req_6186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => addr_of_2532_final_reg_req_1); -- 
    cr_6236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => ptr_deref_2535_store_0_req_1); -- 
    rr_6245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2541_inst_req_0); -- 
    cr_6250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_5730_elements(91), ack => type_cast_2541_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2489_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2519_wire : std_logic_vector(31 downto 0);
    signal R_idxprom102_2530_resized : std_logic_vector(13 downto 0);
    signal R_idxprom102_2530_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2500_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2500_scaled : std_logic_vector(13 downto 0);
    signal add107_2548 : std_logic_vector(31 downto 0);
    signal add49_2472 : std_logic_vector(15 downto 0);
    signal add93_2477 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2501_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2501_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2501_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2501_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2501_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2501_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2531_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2531_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2531_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2531_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2531_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2531_root_address : std_logic_vector(13 downto 0);
    signal arrayidx103_2533 : std_logic_vector(31 downto 0);
    signal arrayidx97_2503 : std_logic_vector(31 downto 0);
    signal call11_2324 : std_logic_vector(15 downto 0);
    signal call13_2327 : std_logic_vector(15 downto 0);
    signal call14_2330 : std_logic_vector(15 downto 0);
    signal call15_2333 : std_logic_vector(15 downto 0);
    signal call17_2336 : std_logic_vector(15 downto 0);
    signal call19_2339 : std_logic_vector(15 downto 0);
    signal call1_2309 : std_logic_vector(15 downto 0);
    signal call3_2312 : std_logic_vector(15 downto 0);
    signal call5_2315 : std_logic_vector(15 downto 0);
    signal call7_2318 : std_logic_vector(15 downto 0);
    signal call9_2321 : std_logic_vector(15 downto 0);
    signal call_2306 : std_logic_vector(15 downto 0);
    signal cmp122_2586 : std_logic_vector(0 downto 0);
    signal cmp137_2611 : std_logic_vector(0 downto 0);
    signal cmp_2555 : std_logic_vector(0 downto 0);
    signal conv100_2512 : std_logic_vector(31 downto 0);
    signal conv106_2542 : std_logic_vector(31 downto 0);
    signal conv110_2356 : std_logic_vector(31 downto 0);
    signal conv118_2581 : std_logic_vector(31 downto 0);
    signal conv121_2360 : std_logic_vector(31 downto 0);
    signal conv133_2606 : std_logic_vector(31 downto 0);
    signal conv136_2364 : std_logic_vector(31 downto 0);
    signal conv96_2482 : std_logic_vector(31 downto 0);
    signal div27_2352 : std_logic_vector(15 downto 0);
    signal div_2346 : std_logic_vector(15 downto 0);
    signal idxprom102_2526 : std_logic_vector(63 downto 0);
    signal idxprom_2496 : std_logic_vector(63 downto 0);
    signal inc126_2596 : std_logic_vector(15 downto 0);
    signal inc_2576 : std_logic_vector(15 downto 0);
    signal indvar_2454 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2568 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2601 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2395 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2389 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2592 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2467 : std_logic_vector(15 downto 0);
    signal ptr_deref_2506_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2506_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2506_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2506_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2506_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2535_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2535_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2535_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr101_2521 : std_logic_vector(31 downto 0);
    signal shr_2491 : std_logic_vector(31 downto 0);
    signal tmp10_2451 : std_logic_vector(15 downto 0);
    signal tmp164_2406 : std_logic_vector(15 downto 0);
    signal tmp165_2411 : std_logic_vector(15 downto 0);
    signal tmp166_2416 : std_logic_vector(15 downto 0);
    signal tmp1_2375 : std_logic_vector(15 downto 0);
    signal tmp2_2421 : std_logic_vector(15 downto 0);
    signal tmp3_2426 : std_logic_vector(15 downto 0);
    signal tmp4_2381 : std_logic_vector(15 downto 0);
    signal tmp5_2386 : std_logic_vector(15 downto 0);
    signal tmp6_2431 : std_logic_vector(15 downto 0);
    signal tmp7_2436 : std_logic_vector(15 downto 0);
    signal tmp8_2441 : std_logic_vector(15 downto 0);
    signal tmp98_2507 : std_logic_vector(63 downto 0);
    signal tmp9_2446 : std_logic_vector(15 downto 0);
    signal tmp_2370 : std_logic_vector(15 downto 0);
    signal type_cast_2344_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2350_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2368_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2379_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2392_wire : std_logic_vector(15 downto 0);
    signal type_cast_2394_wire : std_logic_vector(15 downto 0);
    signal type_cast_2398_wire : std_logic_vector(15 downto 0);
    signal type_cast_2400_wire : std_logic_vector(15 downto 0);
    signal type_cast_2457_wire : std_logic_vector(15 downto 0);
    signal type_cast_2460_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2465_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2480_wire : std_logic_vector(31 downto 0);
    signal type_cast_2485_wire : std_logic_vector(31 downto 0);
    signal type_cast_2488_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2494_wire : std_logic_vector(63 downto 0);
    signal type_cast_2510_wire : std_logic_vector(31 downto 0);
    signal type_cast_2515_wire : std_logic_vector(31 downto 0);
    signal type_cast_2518_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2524_wire : std_logic_vector(63 downto 0);
    signal type_cast_2540_wire : std_logic_vector(31 downto 0);
    signal type_cast_2546_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2551_wire : std_logic_vector(31 downto 0);
    signal type_cast_2553_wire : std_logic_vector(31 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2574_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2579_wire : std_logic_vector(31 downto 0);
    signal type_cast_2604_wire : std_logic_vector(31 downto 0);
    signal type_cast_2622_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2501_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2501_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2501_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2501_resized_base_address <= "00000000000000";
    array_obj_ref_2531_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2531_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2531_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2531_resized_base_address <= "00000000000000";
    ptr_deref_2506_word_offset_0 <= "00000000000000";
    ptr_deref_2535_word_offset_0 <= "00000000000000";
    type_cast_2344_wire_constant <= "0000000000000001";
    type_cast_2350_wire_constant <= "0000000000000001";
    type_cast_2368_wire_constant <= "1111111111111111";
    type_cast_2379_wire_constant <= "1111111111111111";
    type_cast_2460_wire_constant <= "0000000000000000";
    type_cast_2465_wire_constant <= "0000000000000100";
    type_cast_2488_wire_constant <= "00000000000000000000000000000010";
    type_cast_2518_wire_constant <= "00000000000000000000000000000010";
    type_cast_2546_wire_constant <= "00000000000000000000000000000100";
    type_cast_2566_wire_constant <= "0000000000000001";
    type_cast_2574_wire_constant <= "0000000000000001";
    type_cast_2622_wire_constant <= "0000000000000001";
    phi_stmt_2389: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2392_wire & type_cast_2394_wire;
      req <= phi_stmt_2389_req_0 & phi_stmt_2389_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2389",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2389_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2389,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2389
    phi_stmt_2395: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2398_wire & type_cast_2400_wire;
      req <= phi_stmt_2395_req_0 & phi_stmt_2395_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2395",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2395_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2395,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2395
    phi_stmt_2454: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2457_wire & type_cast_2460_wire_constant;
      req <= phi_stmt_2454_req_0 & phi_stmt_2454_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2454",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2454_ack_0,
          idata => idata,
          odata => indvar_2454,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2454
    -- flow-through select operator MUX_2591_inst
    input_dim1x_x2_2592 <= div27_2352 when (cmp122_2586(0) /=  '0') else inc_2576;
    addr_of_2502_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2502_final_reg_req_0;
      addr_of_2502_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2502_final_reg_req_1;
      addr_of_2502_final_reg_ack_1<= rack(0);
      addr_of_2502_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2502_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2501_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx97_2503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2532_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2532_final_reg_req_0;
      addr_of_2532_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2532_final_reg_req_1;
      addr_of_2532_final_reg_ack_1<= rack(0);
      addr_of_2532_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2532_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2531_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx103_2533,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2355_inst_req_0;
      type_cast_2355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2355_inst_req_1;
      type_cast_2355_inst_ack_1<= rack(0);
      type_cast_2355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_2356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2359_inst_req_0;
      type_cast_2359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2359_inst_req_1;
      type_cast_2359_inst_ack_1<= rack(0);
      type_cast_2359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_2309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_2360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2363_inst_req_0;
      type_cast_2363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2363_inst_req_1;
      type_cast_2363_inst_ack_1<= rack(0);
      type_cast_2363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_2364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2392_inst_req_0;
      type_cast_2392_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2392_inst_req_1;
      type_cast_2392_inst_ack_1<= rack(0);
      type_cast_2392_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2392_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2392_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2394_inst_req_0;
      type_cast_2394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2394_inst_req_1;
      type_cast_2394_inst_ack_1<= rack(0);
      type_cast_2394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div27_2352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2394_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2398_inst_req_0;
      type_cast_2398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2398_inst_req_1;
      type_cast_2398_inst_ack_1<= rack(0);
      type_cast_2398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2601,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2398_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2400_inst_req_0;
      type_cast_2400_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2400_inst_req_1;
      type_cast_2400_inst_ack_1<= rack(0);
      type_cast_2400_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2400_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2400_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2457_inst_req_0;
      type_cast_2457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2457_inst_req_1;
      type_cast_2457_inst_ack_1<= rack(0);
      type_cast_2457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2568,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2457_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2481_inst_req_0;
      type_cast_2481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2481_inst_req_1;
      type_cast_2481_inst_ack_1<= rack(0);
      type_cast_2481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2480_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_2482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2485_inst
    process(conv96_2482) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv96_2482(31 downto 0);
      type_cast_2485_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2490_inst
    process(ASHR_i32_i32_2489_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2489_wire(31 downto 0);
      shr_2491 <= tmp_var; -- 
    end process;
    type_cast_2495_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2495_inst_req_0;
      type_cast_2495_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2495_inst_req_1;
      type_cast_2495_inst_ack_1<= rack(0);
      type_cast_2495_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2495_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2494_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2496,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2511_inst_req_0;
      type_cast_2511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2511_inst_req_1;
      type_cast_2511_inst_ack_1<= rack(0);
      type_cast_2511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2510_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_2512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2515_inst
    process(conv100_2512) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv100_2512(31 downto 0);
      type_cast_2515_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2520_inst
    process(ASHR_i32_i32_2519_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2519_wire(31 downto 0);
      shr101_2521 <= tmp_var; -- 
    end process;
    type_cast_2525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2525_inst_req_0;
      type_cast_2525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2525_inst_req_1;
      type_cast_2525_inst_ack_1<= rack(0);
      type_cast_2525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2524_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom102_2526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2541_inst_req_0;
      type_cast_2541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2541_inst_req_1;
      type_cast_2541_inst_ack_1<= rack(0);
      type_cast_2541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2540_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv106_2542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2551_inst
    process(add107_2548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add107_2548(31 downto 0);
      type_cast_2551_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2553_inst
    process(conv110_2356) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv110_2356(31 downto 0);
      type_cast_2553_wire <= tmp_var; -- 
    end process;
    type_cast_2580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2580_inst_req_0;
      type_cast_2580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2580_inst_req_1;
      type_cast_2580_inst_ack_1<= rack(0);
      type_cast_2580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2579_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_2581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2595_inst_req_0;
      type_cast_2595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2595_inst_req_1;
      type_cast_2595_inst_ack_1<= rack(0);
      type_cast_2595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp122_2586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc126_2596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2605_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2605_inst_req_0;
      type_cast_2605_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2605_inst_req_1;
      type_cast_2605_inst_ack_1<= rack(0);
      type_cast_2605_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2605_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2604_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv133_2606,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2501_index_1_rename
    process(R_idxprom_2500_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2500_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2500_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2501_index_1_resize
    process(idxprom_2496) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2496;
      ov := iv(13 downto 0);
      R_idxprom_2500_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2501_root_address_inst
    process(array_obj_ref_2501_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2501_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2501_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2531_index_1_rename
    process(R_idxprom102_2530_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom102_2530_resized;
      ov(13 downto 0) := iv;
      R_idxprom102_2530_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2531_index_1_resize
    process(idxprom102_2526) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom102_2526;
      ov := iv(13 downto 0);
      R_idxprom102_2530_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2531_root_address_inst
    process(array_obj_ref_2531_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2531_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2531_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2506_addr_0
    process(ptr_deref_2506_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2506_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2506_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2506_base_resize
    process(arrayidx97_2503) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx97_2503;
      ov := iv(13 downto 0);
      ptr_deref_2506_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2506_gather_scatter
    process(ptr_deref_2506_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2506_data_0;
      ov(63 downto 0) := iv;
      tmp98_2507 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2506_root_address_inst
    process(ptr_deref_2506_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2506_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2506_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_addr_0
    process(ptr_deref_2535_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2535_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2535_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_base_resize
    process(arrayidx103_2533) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx103_2533;
      ov := iv(13 downto 0);
      ptr_deref_2535_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_gather_scatter
    process(tmp98_2507) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp98_2507;
      ov(63 downto 0) := iv;
      ptr_deref_2535_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2535_root_address_inst
    process(ptr_deref_2535_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2535_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2535_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2556_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2555;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2556_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2556_branch_req_0,
          ack0 => if_stmt_2556_branch_ack_0,
          ack1 => if_stmt_2556_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2612_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp137_2611;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2612_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2612_branch_req_0,
          ack0 => if_stmt_2612_branch_ack_0,
          ack1 => if_stmt_2612_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2369_inst
    process(call9_2321) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2321, type_cast_2368_wire_constant, tmp_var);
      tmp_2370 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2380_inst
    process(call7_2318) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2318, type_cast_2379_wire_constant, tmp_var);
      tmp4_2381 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2410_inst
    process(input_dim1x_x1x_xph_2389, tmp164_2406) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2389, tmp164_2406, tmp_var);
      tmp165_2411 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2425_inst
    process(tmp1_2375, tmp2_2421) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_2375, tmp2_2421, tmp_var);
      tmp3_2426 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2435_inst
    process(tmp5_2386, tmp6_2431) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2386, tmp6_2431, tmp_var);
      tmp7_2436 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2445_inst
    process(tmp3_2426, tmp8_2441) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2426, tmp8_2441, tmp_var);
      tmp9_2446 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2471_inst
    process(tmp166_2416, input_dim2x_x1_2467) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp166_2416, input_dim2x_x1_2467, tmp_var);
      add49_2472 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2476_inst
    process(tmp10_2451, input_dim2x_x1_2467) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2451, input_dim2x_x1_2467, tmp_var);
      add93_2477 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2567_inst
    process(indvar_2454) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2454, type_cast_2566_wire_constant, tmp_var);
      indvarx_xnext_2568 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2575_inst
    process(input_dim1x_x1x_xph_2389) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2389, type_cast_2574_wire_constant, tmp_var);
      inc_2576 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2600_inst
    process(inc126_2596, input_dim0x_x2x_xph_2395) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc126_2596, input_dim0x_x2x_xph_2395, tmp_var);
      input_dim0x_x0_2601 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2547_inst
    process(conv106_2542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv106_2542, type_cast_2546_wire_constant, tmp_var);
      add107_2548 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2489_inst
    process(type_cast_2485_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2485_wire, type_cast_2488_wire_constant, tmp_var);
      ASHR_i32_i32_2489_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2519_inst
    process(type_cast_2515_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2515_wire, type_cast_2518_wire_constant, tmp_var);
      ASHR_i32_i32_2519_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2585_inst
    process(conv118_2581, conv121_2360) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv118_2581, conv121_2360, tmp_var);
      cmp122_2586 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2610_inst
    process(conv133_2606, conv136_2364) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv133_2606, conv136_2364, tmp_var);
      cmp137_2611 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2345_inst
    process(call_2306) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2306, type_cast_2344_wire_constant, tmp_var);
      div_2346 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2351_inst
    process(call1_2309) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call1_2309, type_cast_2350_wire_constant, tmp_var);
      div27_2352 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2405_inst
    process(call1_2309, input_dim0x_x2x_xph_2395) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call1_2309, input_dim0x_x2x_xph_2395, tmp_var);
      tmp164_2406 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2415_inst
    process(call3_2312, tmp165_2411) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call3_2312, tmp165_2411, tmp_var);
      tmp166_2416 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2420_inst
    process(call13_2327, input_dim1x_x1x_xph_2389) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2327, input_dim1x_x1x_xph_2389, tmp_var);
      tmp2_2421 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2430_inst
    process(call13_2327, input_dim0x_x2x_xph_2395) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call13_2327, input_dim0x_x2x_xph_2395, tmp_var);
      tmp6_2431 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2440_inst
    process(call17_2336, tmp7_2436) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call17_2336, tmp7_2436, tmp_var);
      tmp8_2441 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2450_inst
    process(call19_2339, tmp9_2446) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(call19_2339, tmp9_2446, tmp_var);
      tmp10_2451 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2466_inst
    process(indvar_2454) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2454, type_cast_2465_wire_constant, tmp_var);
      input_dim2x_x1_2467 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2554_inst
    process(type_cast_2551_wire, type_cast_2553_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2551_wire, type_cast_2553_wire, tmp_var);
      cmp_2555 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2374_inst
    process(tmp_2370, call14_2330) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_2370, call14_2330, tmp_var);
      tmp1_2375 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2385_inst
    process(tmp4_2381, call14_2330) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2381, call14_2330, tmp_var);
      tmp5_2386 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2501_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2500_scaled;
      array_obj_ref_2501_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2501_index_offset_req_0;
      array_obj_ref_2501_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2501_index_offset_req_1;
      array_obj_ref_2501_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2531_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom102_2530_scaled;
      array_obj_ref_2531_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2531_index_offset_req_0;
      array_obj_ref_2531_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2531_index_offset_req_1;
      array_obj_ref_2531_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_2480_inst
    process(add49_2472) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add49_2472, tmp_var);
      type_cast_2480_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2494_inst
    process(shr_2491) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2491, tmp_var);
      type_cast_2494_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2510_inst
    process(add93_2477) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add93_2477, tmp_var);
      type_cast_2510_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2524_inst
    process(shr101_2521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr101_2521, tmp_var);
      type_cast_2524_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2540_inst
    process(input_dim2x_x1_2467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2467, tmp_var);
      type_cast_2540_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2579_inst
    process(inc_2576) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2576, tmp_var);
      type_cast_2579_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2604_inst
    process(input_dim0x_x0_2601) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2601, tmp_var);
      type_cast_2604_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2506_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2506_load_0_req_0;
      ptr_deref_2506_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2506_load_0_req_1;
      ptr_deref_2506_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2506_word_address_0;
      ptr_deref_2506_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2535_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2535_store_0_req_0;
      ptr_deref_2535_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2535_store_0_req_1;
      ptr_deref_2535_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2535_word_address_0;
      data_in <= ptr_deref_2535_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_2329_inst RPIPE_Block1_start_2332_inst RPIPE_Block1_start_2335_inst RPIPE_Block1_start_2338_inst RPIPE_Block1_start_2326_inst RPIPE_Block1_start_2323_inst RPIPE_Block1_start_2320_inst RPIPE_Block1_start_2317_inst RPIPE_Block1_start_2314_inst RPIPE_Block1_start_2311_inst RPIPE_Block1_start_2308_inst RPIPE_Block1_start_2305_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(191 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_Block1_start_2329_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_2332_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_2335_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_2338_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_2326_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_2323_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_2320_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_2317_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_2314_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_2311_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_2308_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_2305_inst_req_0;
      RPIPE_Block1_start_2329_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_2332_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_2335_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_2338_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_2326_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_2323_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_2320_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_2317_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_2314_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_2311_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_2308_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_2305_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_Block1_start_2329_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_2332_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_2335_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_2338_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_2326_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_2323_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_2320_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_2317_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_2314_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_2311_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_2308_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_2305_inst_req_1;
      RPIPE_Block1_start_2329_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_2332_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_2335_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_2338_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_2326_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_2323_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_2320_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_2317_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_2314_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_2311_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_2308_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_2305_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call14_2330 <= data_out(191 downto 176);
      call15_2333 <= data_out(175 downto 160);
      call17_2336 <= data_out(159 downto 144);
      call19_2339 <= data_out(143 downto 128);
      call13_2327 <= data_out(127 downto 112);
      call11_2324 <= data_out(111 downto 96);
      call9_2321 <= data_out(95 downto 80);
      call7_2318 <= data_out(79 downto 64);
      call5_2315 <= data_out(63 downto 48);
      call3_2312 <= data_out(47 downto 32);
      call1_2309 <= data_out(31 downto 16);
      call_2306 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2620_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2620_inst_req_0;
      WPIPE_Block3_done_2620_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2620_inst_req_1;
      WPIPE_Block3_done_2620_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2622_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_29_load_0_req_0 : boolean;
  signal LOAD_count_29_load_0_ack_0 : boolean;
  signal LOAD_count_29_load_0_req_1 : boolean;
  signal LOAD_count_29_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_30/$entry
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_update_start_
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_30/LOAD_count_29_Sample/$entry
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_29_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_30/LOAD_count_29_Sample/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$entry
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_30/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_30/LOAD_count_29_Update/LOAD_count_29_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_29_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_29_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_29_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_29_word_address_0 <= "0";
    -- equivalence LOAD_count_29_gather_scatter
    process(LOAD_count_29_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_29_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_29_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_29_load_0_req_0;
      LOAD_count_29_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_29_load_0_req_1;
      LOAD_count_29_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_29_word_address_0;
      LOAD_count_29_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Block2_start_pipe_read_data: out std_logic_vector(15 downto 0);
    Block2_start_pipe_read_req : in std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : out std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data: out std_logic_vector(15 downto 0);
    Block3_start_pipe_read_req : in std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(47 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(2 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(2 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(1 downto 1),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(1 downto 1),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(31 downto 16),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(2 downto 2),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(2 downto 2),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(47 downto 32),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 3,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
