-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant input_1_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant input_2_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant output_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  -- 
end package ahir_system_global_package;
