-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_34_start: Boolean;
  signal convTranspose_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block2_start_1081_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_req_0 : boolean;
  signal addr_of_694_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal if_stmt_637_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_1 : boolean;
  signal type_cast_615_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_0 : boolean;
  signal type_cast_615_inst_req_1 : boolean;
  signal type_cast_597_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 : boolean;
  signal type_cast_543_inst_ack_1 : boolean;
  signal type_cast_597_inst_req_0 : boolean;
  signal type_cast_543_inst_req_1 : boolean;
  signal type_cast_543_inst_ack_0 : boolean;
  signal type_cast_543_inst_req_0 : boolean;
  signal array_obj_ref_693_index_offset_req_1 : boolean;
  signal type_cast_1417_inst_ack_0 : boolean;
  signal ptr_deref_623_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_1 : boolean;
  signal ptr_deref_623_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 : boolean;
  signal type_cast_714_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_0 : boolean;
  signal type_cast_44_inst_req_0 : boolean;
  signal type_cast_44_inst_ack_0 : boolean;
  signal type_cast_44_inst_req_1 : boolean;
  signal type_cast_44_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1013_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 : boolean;
  signal type_cast_144_inst_req_0 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal type_cast_144_inst_ack_0 : boolean;
  signal type_cast_714_inst_req_0 : boolean;
  signal type_cast_57_inst_req_0 : boolean;
  signal type_cast_57_inst_ack_0 : boolean;
  signal type_cast_57_inst_req_1 : boolean;
  signal type_cast_57_inst_ack_1 : boolean;
  signal type_cast_664_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_0 : boolean;
  signal type_cast_615_inst_ack_0 : boolean;
  signal array_obj_ref_693_index_offset_ack_0 : boolean;
  signal type_cast_69_inst_req_0 : boolean;
  signal type_cast_69_inst_ack_0 : boolean;
  signal type_cast_69_inst_req_1 : boolean;
  signal type_cast_69_inst_ack_1 : boolean;
  signal type_cast_664_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_0 : boolean;
  signal ptr_deref_623_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 : boolean;
  signal type_cast_1417_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_0 : boolean;
  signal type_cast_615_inst_req_0 : boolean;
  signal array_obj_ref_693_index_offset_req_0 : boolean;
  signal type_cast_82_inst_req_0 : boolean;
  signal ptr_deref_623_store_0_req_0 : boolean;
  signal type_cast_82_inst_ack_0 : boolean;
  signal type_cast_82_inst_req_1 : boolean;
  signal type_cast_82_inst_ack_1 : boolean;
  signal type_cast_664_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_1 : boolean;
  signal type_cast_94_inst_req_0 : boolean;
  signal type_cast_94_inst_ack_0 : boolean;
  signal type_cast_94_inst_req_1 : boolean;
  signal type_cast_94_inst_ack_1 : boolean;
  signal type_cast_714_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_1 : boolean;
  signal type_cast_664_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_req_0 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_1 : boolean;
  signal type_cast_107_inst_req_0 : boolean;
  signal type_cast_107_inst_ack_0 : boolean;
  signal type_cast_107_inst_req_1 : boolean;
  signal type_cast_107_inst_ack_1 : boolean;
  signal type_cast_714_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal type_cast_732_inst_req_1 : boolean;
  signal type_cast_579_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 : boolean;
  signal type_cast_579_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_req_0 : boolean;
  signal type_cast_119_inst_req_0 : boolean;
  signal type_cast_119_inst_ack_0 : boolean;
  signal type_cast_119_inst_req_1 : boolean;
  signal type_cast_119_inst_ack_1 : boolean;
  signal addr_of_694_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal type_cast_132_inst_req_0 : boolean;
  signal type_cast_132_inst_ack_0 : boolean;
  signal type_cast_132_inst_req_1 : boolean;
  signal type_cast_132_inst_ack_1 : boolean;
  signal addr_of_694_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 : boolean;
  signal type_cast_579_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_1 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal type_cast_1387_inst_ack_1 : boolean;
  signal type_cast_144_inst_req_1 : boolean;
  signal type_cast_144_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_0 : boolean;
  signal type_cast_579_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_0 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal type_cast_157_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_0 : boolean;
  signal type_cast_157_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_1 : boolean;
  signal type_cast_732_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 : boolean;
  signal type_cast_169_inst_req_0 : boolean;
  signal type_cast_169_inst_ack_0 : boolean;
  signal type_cast_169_inst_req_1 : boolean;
  signal type_cast_169_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_1 : boolean;
  signal addr_of_694_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_0 : boolean;
  signal type_cast_701_inst_ack_1 : boolean;
  signal type_cast_701_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal ptr_deref_1373_load_0_ack_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal if_stmt_637_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_1 : boolean;
  signal type_cast_207_inst_req_0 : boolean;
  signal type_cast_207_inst_ack_0 : boolean;
  signal type_cast_207_inst_req_1 : boolean;
  signal type_cast_207_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 : boolean;
  signal type_cast_216_inst_req_0 : boolean;
  signal type_cast_216_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_req_0 : boolean;
  signal type_cast_216_inst_req_1 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal type_cast_216_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_1 : boolean;
  signal type_cast_220_inst_req_0 : boolean;
  signal type_cast_220_inst_ack_0 : boolean;
  signal type_cast_220_inst_req_1 : boolean;
  signal type_cast_220_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1016_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_1 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_1 : boolean;
  signal type_cast_261_inst_req_0 : boolean;
  signal type_cast_261_inst_ack_0 : boolean;
  signal type_cast_261_inst_req_1 : boolean;
  signal type_cast_261_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal type_cast_265_inst_req_0 : boolean;
  signal type_cast_265_inst_ack_0 : boolean;
  signal type_cast_265_inst_req_1 : boolean;
  signal type_cast_265_inst_ack_1 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_273_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_0 : boolean;
  signal type_cast_273_inst_req_1 : boolean;
  signal type_cast_273_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 : boolean;
  signal type_cast_701_inst_ack_0 : boolean;
  signal type_cast_701_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_0 : boolean;
  signal type_cast_295_inst_req_0 : boolean;
  signal type_cast_295_inst_ack_0 : boolean;
  signal type_cast_295_inst_req_1 : boolean;
  signal type_cast_295_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_ack_1 : boolean;
  signal type_cast_597_inst_ack_1 : boolean;
  signal type_cast_308_inst_req_0 : boolean;
  signal type_cast_308_inst_ack_0 : boolean;
  signal type_cast_308_inst_req_1 : boolean;
  signal type_cast_308_inst_ack_1 : boolean;
  signal if_stmt_637_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 : boolean;
  signal type_cast_597_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal ptr_deref_1373_load_0_req_1 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 : boolean;
  signal array_obj_ref_693_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_ack_1 : boolean;
  signal type_cast_333_inst_req_0 : boolean;
  signal type_cast_333_inst_ack_0 : boolean;
  signal type_cast_333_inst_req_1 : boolean;
  signal type_cast_333_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal type_cast_1417_inst_req_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 : boolean;
  signal type_cast_1417_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_req_0 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_ack_1 : boolean;
  signal type_cast_383_inst_req_0 : boolean;
  signal type_cast_383_inst_ack_0 : boolean;
  signal type_cast_383_inst_req_1 : boolean;
  signal type_cast_383_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_1 : boolean;
  signal type_cast_395_inst_req_0 : boolean;
  signal type_cast_395_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_1 : boolean;
  signal type_cast_395_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_1 : boolean;
  signal if_stmt_421_branch_req_0 : boolean;
  signal if_stmt_421_branch_ack_1 : boolean;
  signal if_stmt_421_branch_ack_0 : boolean;
  signal if_stmt_436_branch_req_0 : boolean;
  signal if_stmt_436_branch_ack_1 : boolean;
  signal if_stmt_436_branch_ack_0 : boolean;
  signal type_cast_457_inst_req_0 : boolean;
  signal type_cast_457_inst_ack_0 : boolean;
  signal type_cast_457_inst_req_1 : boolean;
  signal type_cast_457_inst_ack_1 : boolean;
  signal array_obj_ref_486_index_offset_req_0 : boolean;
  signal array_obj_ref_486_index_offset_ack_0 : boolean;
  signal array_obj_ref_486_index_offset_req_1 : boolean;
  signal array_obj_ref_486_index_offset_ack_1 : boolean;
  signal addr_of_487_final_reg_req_0 : boolean;
  signal addr_of_487_final_reg_ack_0 : boolean;
  signal addr_of_487_final_reg_req_1 : boolean;
  signal addr_of_487_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_ack_1 : boolean;
  signal type_cast_494_inst_req_0 : boolean;
  signal type_cast_494_inst_ack_0 : boolean;
  signal type_cast_494_inst_req_1 : boolean;
  signal type_cast_494_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_ack_1 : boolean;
  signal type_cast_507_inst_req_0 : boolean;
  signal type_cast_507_inst_ack_0 : boolean;
  signal type_cast_507_inst_req_1 : boolean;
  signal type_cast_507_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_ack_1 : boolean;
  signal type_cast_525_inst_req_0 : boolean;
  signal type_cast_525_inst_ack_0 : boolean;
  signal type_cast_525_inst_req_1 : boolean;
  signal type_cast_525_inst_ack_1 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1013_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1072_inst_ack_1 : boolean;
  signal type_cast_768_inst_req_0 : boolean;
  signal type_cast_768_inst_ack_0 : boolean;
  signal type_cast_768_inst_req_1 : boolean;
  signal type_cast_768_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1013_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_req_1 : boolean;
  signal type_cast_786_inst_req_0 : boolean;
  signal type_cast_786_inst_ack_0 : boolean;
  signal type_cast_786_inst_req_1 : boolean;
  signal type_cast_786_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1013_inst_req_0 : boolean;
  signal type_cast_804_inst_req_0 : boolean;
  signal type_cast_804_inst_ack_0 : boolean;
  signal type_cast_804_inst_req_1 : boolean;
  signal type_cast_804_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_1 : boolean;
  signal type_cast_1387_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1043_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_1 : boolean;
  signal type_cast_822_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_1 : boolean;
  signal type_cast_1061_inst_ack_1 : boolean;
  signal type_cast_1061_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1043_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1072_inst_req_0 : boolean;
  signal ptr_deref_830_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_1 : boolean;
  signal ptr_deref_830_store_0_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_1 : boolean;
  signal WPIPE_Block0_start_999_inst_ack_1 : boolean;
  signal ptr_deref_830_store_0_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_1 : boolean;
  signal ptr_deref_830_store_0_ack_1 : boolean;
  signal if_stmt_844_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_0 : boolean;
  signal if_stmt_844_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_0 : boolean;
  signal if_stmt_844_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_999_inst_req_1 : boolean;
  signal type_cast_855_inst_req_0 : boolean;
  signal type_cast_855_inst_ack_0 : boolean;
  signal type_cast_855_inst_req_1 : boolean;
  signal type_cast_855_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_0 : boolean;
  signal type_cast_1339_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_0 : boolean;
  signal type_cast_859_inst_req_0 : boolean;
  signal type_cast_859_inst_ack_0 : boolean;
  signal type_cast_859_inst_req_1 : boolean;
  signal type_cast_859_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_0 : boolean;
  signal type_cast_1061_inst_ack_0 : boolean;
  signal type_cast_1061_inst_req_0 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1040_inst_ack_1 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal type_cast_863_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1040_inst_req_1 : boolean;
  signal type_cast_863_inst_ack_1 : boolean;
  signal if_stmt_881_branch_req_0 : boolean;
  signal if_stmt_881_branch_ack_1 : boolean;
  signal if_stmt_881_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_1 : boolean;
  signal type_cast_908_inst_req_0 : boolean;
  signal type_cast_908_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_1 : boolean;
  signal type_cast_908_inst_req_1 : boolean;
  signal type_cast_908_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_1 : boolean;
  signal type_cast_1339_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_1 : boolean;
  signal array_obj_ref_937_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1040_inst_ack_0 : boolean;
  signal array_obj_ref_937_index_offset_ack_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal array_obj_ref_937_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1040_inst_req_0 : boolean;
  signal array_obj_ref_937_index_offset_ack_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_1 : boolean;
  signal addr_of_938_final_reg_req_0 : boolean;
  signal addr_of_938_final_reg_ack_0 : boolean;
  signal addr_of_938_final_reg_req_1 : boolean;
  signal addr_of_938_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_1 : boolean;
  signal WPIPE_Block0_start_999_inst_ack_0 : boolean;
  signal ptr_deref_941_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_0 : boolean;
  signal ptr_deref_941_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_0 : boolean;
  signal WPIPE_Block0_start_999_inst_req_0 : boolean;
  signal ptr_deref_941_store_0_req_1 : boolean;
  signal ptr_deref_941_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_1 : boolean;
  signal if_stmt_956_branch_req_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_1 : boolean;
  signal if_stmt_956_branch_ack_1 : boolean;
  signal if_stmt_956_branch_ack_0 : boolean;
  signal call_stmt_967_call_req_0 : boolean;
  signal call_stmt_967_call_ack_0 : boolean;
  signal WPIPE_Block1_start_1069_inst_ack_1 : boolean;
  signal call_stmt_967_call_req_1 : boolean;
  signal call_stmt_967_call_ack_1 : boolean;
  signal type_cast_1397_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_0 : boolean;
  signal type_cast_972_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_0 : boolean;
  signal type_cast_972_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1069_inst_req_1 : boolean;
  signal type_cast_972_inst_req_1 : boolean;
  signal type_cast_972_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_req_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_1 : boolean;
  signal type_cast_1387_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1096_inst_req_0 : boolean;
  signal ptr_deref_1373_load_0_ack_0 : boolean;
  signal WPIPE_Block2_start_1096_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1096_inst_req_1 : boolean;
  signal ptr_deref_1373_load_0_req_0 : boolean;
  signal WPIPE_Block2_start_1096_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_req_1 : boolean;
  signal type_cast_1339_inst_ack_0 : boolean;
  signal type_cast_1387_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1099_inst_ack_1 : boolean;
  signal type_cast_1339_inst_req_0 : boolean;
  signal type_cast_1427_inst_ack_1 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1427_inst_req_1 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal type_cast_1407_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1112_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1112_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1299_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1112_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1112_inst_ack_1 : boolean;
  signal type_cast_1117_inst_req_0 : boolean;
  signal type_cast_1117_inst_ack_0 : boolean;
  signal type_cast_1117_inst_req_1 : boolean;
  signal type_cast_1117_inst_ack_1 : boolean;
  signal type_cast_1377_inst_ack_1 : boolean;
  signal type_cast_1377_inst_req_1 : boolean;
  signal type_cast_1407_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1452_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1455_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0 : boolean;
  signal type_cast_1427_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_1 : boolean;
  signal type_cast_1377_inst_ack_0 : boolean;
  signal type_cast_1407_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1458_inst_req_0 : boolean;
  signal type_cast_1377_inst_req_0 : boolean;
  signal type_cast_1407_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_1 : boolean;
  signal if_stmt_1312_branch_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1296_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1449_inst_req_0 : boolean;
  signal if_stmt_1312_branch_ack_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_1 : boolean;
  signal addr_of_1369_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_1 : boolean;
  signal type_cast_1427_inst_req_0 : boolean;
  signal if_stmt_1312_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_0 : boolean;
  signal addr_of_1369_final_reg_req_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1152_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_req_1 : boolean;
  signal addr_of_1369_final_reg_ack_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_ack_1 : boolean;
  signal type_cast_1447_inst_ack_1 : boolean;
  signal type_cast_1447_inst_req_1 : boolean;
  signal type_cast_1397_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_req_0 : boolean;
  signal addr_of_1369_final_reg_req_0 : boolean;
  signal WPIPE_Block3_start_1155_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1155_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 : boolean;
  signal type_cast_1447_inst_ack_0 : boolean;
  signal type_cast_1447_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_req_1 : boolean;
  signal type_cast_1166_inst_req_0 : boolean;
  signal type_cast_1166_inst_ack_0 : boolean;
  signal type_cast_1166_inst_req_1 : boolean;
  signal type_cast_1166_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_ack_0 : boolean;
  signal type_cast_1397_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1168_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1168_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1168_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1168_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1308_inst_req_0 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal array_obj_ref_1368_index_offset_ack_1 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1293_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_0 : boolean;
  signal array_obj_ref_1368_index_offset_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_1 : boolean;
  signal array_obj_ref_1368_index_offset_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_1 : boolean;
  signal type_cast_1437_inst_ack_1 : boolean;
  signal type_cast_1437_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_0 : boolean;
  signal array_obj_ref_1368_index_offset_req_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_1 : boolean;
  signal type_cast_1437_inst_ack_0 : boolean;
  signal type_cast_1437_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1305_inst_req_0 : boolean;
  signal type_cast_1397_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1290_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1189_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1189_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1189_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1189_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1192_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1192_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1192_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1192_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1195_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1195_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1195_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1195_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1198_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1198_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1198_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1198_inst_ack_1 : boolean;
  signal call_stmt_1202_call_req_0 : boolean;
  signal call_stmt_1202_call_ack_0 : boolean;
  signal call_stmt_1202_call_req_1 : boolean;
  signal call_stmt_1202_call_ack_1 : boolean;
  signal type_cast_1206_inst_req_0 : boolean;
  signal type_cast_1206_inst_ack_0 : boolean;
  signal type_cast_1206_inst_req_1 : boolean;
  signal type_cast_1206_inst_ack_1 : boolean;
  signal type_cast_1215_inst_req_0 : boolean;
  signal type_cast_1215_inst_ack_0 : boolean;
  signal type_cast_1215_inst_req_1 : boolean;
  signal type_cast_1215_inst_ack_1 : boolean;
  signal type_cast_1225_inst_req_0 : boolean;
  signal type_cast_1225_inst_ack_0 : boolean;
  signal type_cast_1225_inst_req_1 : boolean;
  signal type_cast_1225_inst_ack_1 : boolean;
  signal type_cast_1235_inst_req_0 : boolean;
  signal type_cast_1235_inst_ack_0 : boolean;
  signal type_cast_1235_inst_req_1 : boolean;
  signal type_cast_1235_inst_ack_1 : boolean;
  signal type_cast_1245_inst_req_0 : boolean;
  signal type_cast_1245_inst_ack_0 : boolean;
  signal type_cast_1245_inst_req_1 : boolean;
  signal type_cast_1245_inst_ack_1 : boolean;
  signal type_cast_1255_inst_req_0 : boolean;
  signal type_cast_1255_inst_ack_0 : boolean;
  signal type_cast_1255_inst_req_1 : boolean;
  signal type_cast_1255_inst_ack_1 : boolean;
  signal type_cast_1265_inst_req_0 : boolean;
  signal type_cast_1265_inst_ack_0 : boolean;
  signal type_cast_1265_inst_req_1 : boolean;
  signal type_cast_1265_inst_ack_1 : boolean;
  signal type_cast_1275_inst_req_0 : boolean;
  signal type_cast_1275_inst_ack_0 : boolean;
  signal type_cast_1275_inst_req_1 : boolean;
  signal type_cast_1275_inst_ack_1 : boolean;
  signal type_cast_1285_inst_req_0 : boolean;
  signal type_cast_1285_inst_ack_0 : boolean;
  signal type_cast_1285_inst_req_1 : boolean;
  signal type_cast_1285_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1467_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1470_inst_ack_1 : boolean;
  signal if_stmt_1484_branch_req_0 : boolean;
  signal if_stmt_1484_branch_ack_1 : boolean;
  signal if_stmt_1484_branch_ack_0 : boolean;
  signal phi_stmt_474_req_0 : boolean;
  signal type_cast_480_inst_req_0 : boolean;
  signal type_cast_480_inst_ack_0 : boolean;
  signal type_cast_480_inst_req_1 : boolean;
  signal type_cast_480_inst_ack_1 : boolean;
  signal phi_stmt_474_req_1 : boolean;
  signal phi_stmt_474_ack_0 : boolean;
  signal phi_stmt_681_req_0 : boolean;
  signal type_cast_687_inst_req_0 : boolean;
  signal type_cast_687_inst_ack_0 : boolean;
  signal type_cast_687_inst_req_1 : boolean;
  signal type_cast_687_inst_ack_1 : boolean;
  signal phi_stmt_681_req_1 : boolean;
  signal phi_stmt_681_ack_0 : boolean;
  signal phi_stmt_925_req_1 : boolean;
  signal type_cast_928_inst_req_0 : boolean;
  signal type_cast_928_inst_ack_0 : boolean;
  signal type_cast_928_inst_req_1 : boolean;
  signal type_cast_928_inst_ack_1 : boolean;
  signal phi_stmt_925_req_0 : boolean;
  signal phi_stmt_925_ack_0 : boolean;
  signal phi_stmt_1356_req_0 : boolean;
  signal type_cast_1362_inst_req_0 : boolean;
  signal type_cast_1362_inst_ack_0 : boolean;
  signal type_cast_1362_inst_req_1 : boolean;
  signal type_cast_1362_inst_ack_1 : boolean;
  signal phi_stmt_1356_req_1 : boolean;
  signal phi_stmt_1356_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_34: Block -- control-path 
    signal convTranspose_CP_34_elements: BooleanArray(497 downto 0);
    -- 
  begin -- 
    convTranspose_CP_34_elements(0) <= convTranspose_CP_34_start;
    convTranspose_CP_34_symbol <= convTranspose_CP_34_elements(497);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_38/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/branch_block_stmt_38__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/cr
      -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_0); -- 
    cr_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_44_inst_req_1); -- 
    cr_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_57_inst_req_1); -- 
    cr_207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_69_inst_req_1); -- 
    cr_235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_82_inst_req_1); -- 
    cr_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_94_inst_req_1); -- 
    cr_291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_107_inst_req_1); -- 
    cr_319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_119_inst_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_132_inst_req_1); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_345_inst_req_1); -- 
    cr_375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_144_inst_req_1); -- 
    cr_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_157_inst_req_1); -- 
    cr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_169_inst_req_1); -- 
    cr_459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_182_inst_req_1); -- 
    cr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_194_inst_req_1); -- 
    cr_515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_207_inst_req_1); -- 
    cr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_216_inst_req_1); -- 
    cr_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_220_inst_req_1); -- 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_224_inst_req_1); -- 
    cr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_261_inst_req_1); -- 
    cr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_265_inst_req_1); -- 
    cr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_269_inst_req_1); -- 
    cr_613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_273_inst_req_1); -- 
    cr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_295_inst_req_1); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_308_inst_req_1); -- 
    cr_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_320_inst_req_1); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_333_inst_req_1); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_358_inst_req_1); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_370_inst_req_1); -- 
    cr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_383_inst_req_1); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_395_inst_req_1); -- 
    cr_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_408_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_update_start_
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/cr
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_0, ack => convTranspose_CP_34_elements(1)); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(1), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_sample_start_
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_1, ack => convTranspose_CP_34_elements(2)); -- 
    rr_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => type_cast_44_inst_req_0); -- 
    rr_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/ra
      -- 
    ra_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_0, ack => convTranspose_CP_34_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/ca
      -- 
    ca_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_1, ack => convTranspose_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_update_start_
      -- 
    ra_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_0, ack => convTranspose_CP_34_elements(5)); -- 
    cr_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(5), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/rr
      -- 
    ca_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_1, ack => convTranspose_CP_34_elements(6)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => type_cast_57_inst_req_0); -- 
    rr_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_0, ack => convTranspose_CP_34_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/ca
      -- 
    ca_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_1, ack => convTranspose_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_update_start_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/cr
      -- 
    ra_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_0, ack => convTranspose_CP_34_elements(9)); -- 
    cr_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(9), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/rr
      -- 
    ca_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_1, ack => convTranspose_CP_34_elements(10)); -- 
    rr_202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => type_cast_69_inst_req_0); -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/ra
      -- 
    ra_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_0, ack => convTranspose_CP_34_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/ca
      -- 
    ca_208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_1, ack => convTranspose_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_update_start_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/cr
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_0, ack => convTranspose_CP_34_elements(13)); -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(13), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/rr
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_1, ack => convTranspose_CP_34_elements(14)); -- 
    rr_230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => type_cast_82_inst_req_0); -- 
    rr_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/ra
      -- 
    ra_231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_0, ack => convTranspose_CP_34_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/ca
      -- 
    ca_236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_1, ack => convTranspose_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_update_start_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/cr
      -- 
    ra_245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_0, ack => convTranspose_CP_34_elements(17)); -- 
    cr_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(17), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/rr
      -- 
    ca_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_1, ack => convTranspose_CP_34_elements(18)); -- 
    rr_258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => type_cast_94_inst_req_0); -- 
    rr_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/ra
      -- 
    ra_259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_0, ack => convTranspose_CP_34_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/ca
      -- 
    ca_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_1, ack => convTranspose_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_update_start_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/cr
      -- 
    ra_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_0, ack => convTranspose_CP_34_elements(21)); -- 
    cr_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(21), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/rr
      -- 
    ca_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_1, ack => convTranspose_CP_34_elements(22)); -- 
    rr_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => type_cast_107_inst_req_0); -- 
    rr_300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/ra
      -- 
    ra_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_0, ack => convTranspose_CP_34_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/ca
      -- 
    ca_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_1, ack => convTranspose_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_update_start_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/cr
      -- 
    ra_301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_0, ack => convTranspose_CP_34_elements(25)); -- 
    cr_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(25), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/rr
      -- 
    ca_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_1, ack => convTranspose_CP_34_elements(26)); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => type_cast_119_inst_req_0); -- 
    rr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_0, ack => convTranspose_CP_34_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/ca
      -- 
    ca_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_1, ack => convTranspose_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_update_start_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/cr
      -- 
    ra_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_0, ack => convTranspose_CP_34_elements(29)); -- 
    cr_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(29), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/rr
      -- 
    ca_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_1, ack => convTranspose_CP_34_elements(30)); -- 
    rr_342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => type_cast_132_inst_req_0); -- 
    rr_356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/ra
      -- 
    ra_343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_0, ack => convTranspose_CP_34_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_1, ack => convTranspose_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_update_start_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/cr
      -- 
    ra_357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_0, ack => convTranspose_CP_34_elements(33)); -- 
    cr_361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(33), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/rr
      -- 
    ca_362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_1, ack => convTranspose_CP_34_elements(34)); -- 
    rr_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_0); -- 
    rr_370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => type_cast_144_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/ra
      -- 
    ra_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_0, ack => convTranspose_CP_34_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/ca
      -- 
    ca_376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_1, ack => convTranspose_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_update_start_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/cr
      -- 
    ra_385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_0, ack => convTranspose_CP_34_elements(37)); -- 
    cr_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(37), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/rr
      -- 
    ca_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_1, ack => convTranspose_CP_34_elements(38)); -- 
    rr_398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => type_cast_157_inst_req_0); -- 
    rr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/ra
      -- 
    ra_399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_0, ack => convTranspose_CP_34_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/ca
      -- 
    ca_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_1, ack => convTranspose_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_update_start_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/cr
      -- 
    ra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_0, ack => convTranspose_CP_34_elements(41)); -- 
    cr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(41), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/rr
      -- 
    ca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_1, ack => convTranspose_CP_34_elements(42)); -- 
    rr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => type_cast_169_inst_req_0); -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/ra
      -- 
    ra_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_0, ack => convTranspose_CP_34_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/ca
      -- 
    ca_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_1, ack => convTranspose_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_update_start_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/cr
      -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_0, ack => convTranspose_CP_34_elements(45)); -- 
    cr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(45), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/rr
      -- 
    ca_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_1, ack => convTranspose_CP_34_elements(46)); -- 
    rr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_0); -- 
    rr_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => type_cast_182_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/ra
      -- 
    ra_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => convTranspose_CP_34_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/ca
      -- 
    ca_460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => convTranspose_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_update_start_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/cr
      -- 
    ra_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_0, ack => convTranspose_CP_34_elements(49)); -- 
    cr_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(49), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/rr
      -- 
    ca_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_1, ack => convTranspose_CP_34_elements(50)); -- 
    rr_496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_0); -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => type_cast_194_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/ra
      -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => convTranspose_CP_34_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/ca
      -- 
    ca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => convTranspose_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_update_start_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/cr
      -- 
    ra_497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_0, ack => convTranspose_CP_34_elements(53)); -- 
    cr_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(53), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/rr
      -- 
    ca_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_1, ack => convTranspose_CP_34_elements(54)); -- 
    rr_510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => type_cast_207_inst_req_0); -- 
    rr_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/ra
      -- 
    ra_511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_0, ack => convTranspose_CP_34_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/ca
      -- 
    ca_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_1, ack => convTranspose_CP_34_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/rr
      -- 
    rr_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(57), ack => type_cast_216_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(4) & convTranspose_CP_34_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/ra
      -- 
    ra_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_216_inst_ack_0, ack => convTranspose_CP_34_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/ca
      -- 
    ca_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_216_inst_ack_1, ack => convTranspose_CP_34_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/rr
      -- 
    rr_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(60), ack => type_cast_220_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(12) & convTranspose_CP_34_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/ra
      -- 
    ra_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_0, ack => convTranspose_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/ca
      -- 
    ca_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_1, ack => convTranspose_CP_34_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/rr
      -- 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(63), ack => type_cast_224_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(20) & convTranspose_CP_34_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/ra
      -- 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_0, ack => convTranspose_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/ca
      -- 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_1, ack => convTranspose_CP_34_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	28 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/rr
      -- 
    rr_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(66), ack => type_cast_261_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(32) & convTranspose_CP_34_elements(28);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/ra
      -- 
    ra_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_0, ack => convTranspose_CP_34_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/ca
      -- 
    ca_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_1, ack => convTranspose_CP_34_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	36 
    -- CP-element group 69: 	40 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/rr
      -- 
    rr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(69), ack => type_cast_265_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(36) & convTranspose_CP_34_elements(40);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/ra
      -- 
    ra_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_0, ack => convTranspose_CP_34_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/ca
      -- 
    ca_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_1, ack => convTranspose_CP_34_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/rr
      -- 
    rr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(72), ack => type_cast_269_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(44) & convTranspose_CP_34_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/ra
      -- 
    ra_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => convTranspose_CP_34_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/ca
      -- 
    ca_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => convTranspose_CP_34_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/rr
      -- 
    rr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(75), ack => type_cast_273_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(52) & convTranspose_CP_34_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/ra
      -- 
    ra_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_0, ack => convTranspose_CP_34_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/ca
      -- 
    ca_614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_1, ack => convTranspose_CP_34_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_update_start_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/cr
      -- 
    ra_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_0, ack => convTranspose_CP_34_elements(78)); -- 
    cr_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(78), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/rr
      -- 
    ca_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_1, ack => convTranspose_CP_34_elements(79)); -- 
    rr_636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => type_cast_295_inst_req_0); -- 
    rr_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => RPIPE_ConvTranspose_input_pipe_304_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/ra
      -- 
    ra_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_0, ack => convTranspose_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/ca
      -- 
    ca_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_1, ack => convTranspose_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_update_start_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/cr
      -- 
    ra_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_304_inst_ack_0, ack => convTranspose_CP_34_elements(82)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(82), ack => RPIPE_ConvTranspose_input_pipe_304_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/rr
      -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_304_inst_ack_1, ack => convTranspose_CP_34_elements(83)); -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => type_cast_308_inst_req_0); -- 
    rr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/ra
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_308_inst_ack_0, ack => convTranspose_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_308_inst_ack_1, ack => convTranspose_CP_34_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_update_start_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/cr
      -- 
    ra_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_0, ack => convTranspose_CP_34_elements(86)); -- 
    cr_683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(86), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/rr
      -- 
    ca_684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_1, ack => convTranspose_CP_34_elements(87)); -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => type_cast_320_inst_req_0); -- 
    rr_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => convTranspose_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/ca
      -- 
    ca_698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => convTranspose_CP_34_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_update_start_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/cr
      -- 
    ra_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_0, ack => convTranspose_CP_34_elements(90)); -- 
    cr_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(90), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/rr
      -- 
    ca_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_1, ack => convTranspose_CP_34_elements(91)); -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => type_cast_333_inst_req_0); -- 
    rr_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/ra
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_0, ack => convTranspose_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/ca
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_1, ack => convTranspose_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_update_start_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/cr
      -- 
    ra_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_0, ack => convTranspose_CP_34_elements(94)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(94), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/rr
      -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_1, ack => convTranspose_CP_34_elements(95)); -- 
    rr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => type_cast_345_inst_req_0); -- 
    rr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/ra
      -- 
    ra_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => convTranspose_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_update_completed_
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => convTranspose_CP_34_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_update_start_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/cr
      -- 
    ra_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_0, ack => convTranspose_CP_34_elements(98)); -- 
    cr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(98), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/rr
      -- 
    ca_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_1, ack => convTranspose_CP_34_elements(99)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => type_cast_358_inst_req_0); -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/ra
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => convTranspose_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/ca
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => convTranspose_CP_34_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_update_start_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/cr
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_0, ack => convTranspose_CP_34_elements(102)); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(102), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/rr
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_1, ack => convTranspose_CP_34_elements(103)); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => type_cast_370_inst_req_0); -- 
    rr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => RPIPE_ConvTranspose_input_pipe_379_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/ra
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => convTranspose_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/ca
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => convTranspose_CP_34_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_update_start_
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/cr
      -- 
    ra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_379_inst_ack_0, ack => convTranspose_CP_34_elements(106)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(106), ack => RPIPE_ConvTranspose_input_pipe_379_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/rr
      -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_379_inst_ack_1, ack => convTranspose_CP_34_elements(107)); -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => type_cast_383_inst_req_0); -- 
    rr_846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/ra
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_0, ack => convTranspose_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/ca
      -- 
    ca_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_1, ack => convTranspose_CP_34_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_update_start_
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/cr
      -- 
    ra_847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_0, ack => convTranspose_CP_34_elements(110)); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(110), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/rr
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_1, ack => convTranspose_CP_34_elements(111)); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => type_cast_395_inst_req_0); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => RPIPE_ConvTranspose_input_pipe_404_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/ra
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_0, ack => convTranspose_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/ca
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_1, ack => convTranspose_CP_34_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_update_start_
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/cr
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_404_inst_ack_0, ack => convTranspose_CP_34_elements(114)); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(114), ack => RPIPE_ConvTranspose_input_pipe_404_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/rr
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_404_inst_ack_1, ack => convTranspose_CP_34_elements(115)); -- 
    rr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(115), ack => type_cast_408_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/ra
      -- 
    ra_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_0, ack => convTranspose_CP_34_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/ca
      -- 
    ca_894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_1, ack => convTranspose_CP_34_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420__exit__
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421__entry__
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_38/R_cmp513_422_place
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_else_link/$entry
      -- 
    branch_req_902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(118), ack => if_stmt_421_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(65) & convTranspose_CP_34_elements(62) & convTranspose_CP_34_elements(59) & convTranspose_CP_34_elements(68) & convTranspose_CP_34_elements(77) & convTranspose_CP_34_elements(81) & convTranspose_CP_34_elements(85) & convTranspose_CP_34_elements(89) & convTranspose_CP_34_elements(71) & convTranspose_CP_34_elements(74) & convTranspose_CP_34_elements(93) & convTranspose_CP_34_elements(97) & convTranspose_CP_34_elements(101) & convTranspose_CP_34_elements(105) & convTranspose_CP_34_elements(109) & convTranspose_CP_34_elements(113) & convTranspose_CP_34_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442__exit__
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471__entry__
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_421_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_421_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_update_start_
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/dummy
      -- 
    if_choice_transition_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_421_branch_ack_1, ack => convTranspose_CP_34_elements(119)); -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_457_inst_req_0); -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_457_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	470 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_421_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_421_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_421_branch_ack_0, ack => convTranspose_CP_34_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	470 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643__exit__
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678__entry__
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_update_start_
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_436_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_436_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/dummy
      -- 
    if_choice_transition_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_1, ack => convTranspose_CP_34_elements(121)); -- 
    cr_1310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_664_inst_req_1); -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_664_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	470 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	483 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_38/if_stmt_436_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_38/if_stmt_436_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_0, ack => convTranspose_CP_34_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/ra
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_0, ack => convTranspose_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	471 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471__exit__
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/$exit
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/$entry
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$entry
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_1, ack => convTranspose_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	476 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/ack
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_486_index_offset_ack_0, ack => convTranspose_CP_34_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	476 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/req
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_486_index_offset_ack_1, ack => convTranspose_CP_34_elements(126)); -- 
    req_995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(126), ack => addr_of_487_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/ack
      -- 
    ack_996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_487_final_reg_ack_0, ack => convTranspose_CP_34_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	476 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/ack
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_487_final_reg_ack_1, ack => convTranspose_CP_34_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	476 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_update_start_
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/cr
      -- 
    ra_1010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_490_inst_ack_0, ack => convTranspose_CP_34_elements(129)); -- 
    cr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(129), ack => RPIPE_ConvTranspose_input_pipe_490_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/rr
      -- 
    ca_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_490_inst_ack_1, ack => convTranspose_CP_34_elements(130)); -- 
    rr_1023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => type_cast_494_inst_req_0); -- 
    rr_1037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => RPIPE_ConvTranspose_input_pipe_503_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/ra
      -- 
    ra_1024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_0, ack => convTranspose_CP_34_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	476 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/ca
      -- 
    ca_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_1, ack => convTranspose_CP_34_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_update_start_
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/cr
      -- 
    ra_1038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_503_inst_ack_0, ack => convTranspose_CP_34_elements(133)); -- 
    cr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(133), ack => RPIPE_ConvTranspose_input_pipe_503_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/rr
      -- 
    ca_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_503_inst_ack_1, ack => convTranspose_CP_34_elements(134)); -- 
    rr_1051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => type_cast_507_inst_req_0); -- 
    rr_1065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => RPIPE_ConvTranspose_input_pipe_521_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/ra
      -- 
    ra_1052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_0, ack => convTranspose_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	476 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/ca
      -- 
    ca_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_1, ack => convTranspose_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_update_start_
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/cr
      -- 
    ra_1066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_521_inst_ack_0, ack => convTranspose_CP_34_elements(137)); -- 
    cr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(137), ack => RPIPE_ConvTranspose_input_pipe_521_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/rr
      -- 
    ca_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_521_inst_ack_1, ack => convTranspose_CP_34_elements(138)); -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => type_cast_525_inst_req_0); -- 
    rr_1093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => RPIPE_ConvTranspose_input_pipe_539_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_0, ack => convTranspose_CP_34_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	476 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/ca
      -- 
    ca_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_1, ack => convTranspose_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_update_start_
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_sample_completed_
      -- 
    ra_1094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_539_inst_ack_0, ack => convTranspose_CP_34_elements(141)); -- 
    cr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(141), ack => RPIPE_ConvTranspose_input_pipe_539_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/ca
      -- 
    ca_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_539_inst_ack_1, ack => convTranspose_CP_34_elements(142)); -- 
    rr_1107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => type_cast_543_inst_req_0); -- 
    rr_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_sample_completed_
      -- 
    ra_1108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_0, ack => convTranspose_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	476 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_update_completed_
      -- 
    ca_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_1, ack => convTranspose_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_update_start_
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/$exit
      -- 
    ra_1122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_0, ack => convTranspose_CP_34_elements(145)); -- 
    cr_1126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(145), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/$exit
      -- 
    ca_1127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_1, ack => convTranspose_CP_34_elements(146)); -- 
    rr_1135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => type_cast_561_inst_req_0); -- 
    rr_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => RPIPE_ConvTranspose_input_pipe_575_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_sample_completed_
      -- 
    ra_1136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => convTranspose_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	476 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_update_completed_
      -- 
    ca_1141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => convTranspose_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_update_start_
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_sample_completed_
      -- 
    ra_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_575_inst_ack_0, ack => convTranspose_CP_34_elements(149)); -- 
    cr_1154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(149), ack => RPIPE_ConvTranspose_input_pipe_575_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_update_completed_
      -- 
    ca_1155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_575_inst_ack_1, ack => convTranspose_CP_34_elements(150)); -- 
    rr_1163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => type_cast_579_inst_req_0); -- 
    rr_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_sample_completed_
      -- 
    ra_1164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_0, ack => convTranspose_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	476 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_update_completed_
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_1, ack => convTranspose_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_update_start_
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_sample_completed_
      -- 
    ra_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_0, ack => convTranspose_CP_34_elements(153)); -- 
    cr_1182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(153), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_sample_start_
      -- 
    ca_1183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_1, ack => convTranspose_CP_34_elements(154)); -- 
    rr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => type_cast_597_inst_req_0); -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/$exit
      -- 
    ra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_0, ack => convTranspose_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	476 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/$exit
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_1, ack => convTranspose_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_update_start_
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_sample_completed_
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_0, ack => convTranspose_CP_34_elements(157)); -- 
    cr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(157), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_update_completed_
      -- 
    ca_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_1, ack => convTranspose_CP_34_elements(158)); -- 
    rr_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(158), ack => type_cast_615_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_sample_completed_
      -- 
    ra_1220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_0, ack => convTranspose_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	476 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_update_completed_
      -- 
    ca_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_1, ack => convTranspose_CP_34_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_sample_start_
      -- 
    rr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(161), ack => ptr_deref_623_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(128) & convTranspose_CP_34_elements(132) & convTranspose_CP_34_elements(136) & convTranspose_CP_34_elements(140) & convTranspose_CP_34_elements(144) & convTranspose_CP_34_elements(148) & convTranspose_CP_34_elements(152) & convTranspose_CP_34_elements(156) & convTranspose_CP_34_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_sample_completed_
      -- 
    ra_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_623_store_0_ack_0, ack => convTranspose_CP_34_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	476 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_update_completed_
      -- 
    ca_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_623_store_0_ack_1, ack => convTranspose_CP_34_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	125 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636__exit__
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637__entry__
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/R_exitcond3_638_place
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/$exit
      -- 
    branch_req_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(164), ack => if_stmt_637_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(125) & convTranspose_CP_34_elements(163);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	470 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427__exit__
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_38/if_stmt_637_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_38/if_stmt_637_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_637_branch_ack_1, ack => convTranspose_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	472 
    -- CP-element group 166: 	473 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_38/if_stmt_637_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_38/if_stmt_637_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_637_branch_ack_0, ack => convTranspose_CP_34_elements(166)); -- 
    rr_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_480_inst_req_0); -- 
    cr_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_480_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_sample_completed_
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_0, ack => convTranspose_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	477 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678__exit__
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/$exit
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/$entry
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$entry
      -- 
    ca_1311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_1, ack => convTranspose_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	482 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_sample_complete
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_693_index_offset_ack_0, ack => convTranspose_CP_34_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	482 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/req
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/ack
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_693_index_offset_ack_1, ack => convTranspose_CP_34_elements(170)); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(170), ack => addr_of_694_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/ack
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_694_final_reg_ack_0, ack => convTranspose_CP_34_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	482 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/root_register_ack
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_694_final_reg_ack_1, ack => convTranspose_CP_34_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	482 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_update_start_
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_sample_completed_
      -- 
    ra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_697_inst_ack_0, ack => convTranspose_CP_34_elements(173)); -- 
    cr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(173), ack => RPIPE_ConvTranspose_input_pipe_697_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/$entry
      -- 
    ca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_697_inst_ack_1, ack => convTranspose_CP_34_elements(174)); -- 
    rr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => type_cast_701_inst_req_0); -- 
    rr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => RPIPE_ConvTranspose_input_pipe_710_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/$exit
      -- 
    ra_1383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_0, ack => convTranspose_CP_34_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	482 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_update_completed_
      -- 
    ca_1388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_1, ack => convTranspose_CP_34_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_update_start_
      -- 
    ra_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_710_inst_ack_0, ack => convTranspose_CP_34_elements(177)); -- 
    cr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(177), ack => RPIPE_ConvTranspose_input_pipe_710_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/$entry
      -- 
    ca_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_710_inst_ack_1, ack => convTranspose_CP_34_elements(178)); -- 
    rr_1410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => type_cast_714_inst_req_0); -- 
    rr_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_sample_completed_
      -- 
    ra_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_0, ack => convTranspose_CP_34_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	482 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_update_completed_
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_1, ack => convTranspose_CP_34_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_update_start_
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/$exit
      -- 
    ra_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_0, ack => convTranspose_CP_34_elements(181)); -- 
    cr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(181), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_update_completed_
      -- 
    ca_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_1, ack => convTranspose_CP_34_elements(182)); -- 
    rr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => type_cast_732_inst_req_0); -- 
    rr_1452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => RPIPE_ConvTranspose_input_pipe_746_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/ra
      -- 
    ra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_0, ack => convTranspose_CP_34_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	482 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/$exit
      -- 
    ca_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_1, ack => convTranspose_CP_34_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_update_start_
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_sample_completed_
      -- 
    ra_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_746_inst_ack_0, ack => convTranspose_CP_34_elements(185)); -- 
    cr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(185), ack => RPIPE_ConvTranspose_input_pipe_746_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/rr
      -- 
    ca_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_746_inst_ack_1, ack => convTranspose_CP_34_elements(186)); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => type_cast_750_inst_req_0); -- 
    rr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => RPIPE_ConvTranspose_input_pipe_764_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/ra
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => convTranspose_CP_34_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	482 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/ca
      -- 
    ca_1472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => convTranspose_CP_34_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_update_start_
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/cr
      -- 
    ra_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_764_inst_ack_0, ack => convTranspose_CP_34_elements(189)); -- 
    cr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(189), ack => RPIPE_ConvTranspose_input_pipe_764_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/rr
      -- 
    ca_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_764_inst_ack_1, ack => convTranspose_CP_34_elements(190)); -- 
    rr_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => type_cast_768_inst_req_0); -- 
    rr_1508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => RPIPE_ConvTranspose_input_pipe_782_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/ra
      -- 
    ra_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_0, ack => convTranspose_CP_34_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	482 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/ca
      -- 
    ca_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_1, ack => convTranspose_CP_34_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_update_start_
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/cr
      -- 
    ra_1509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_782_inst_ack_0, ack => convTranspose_CP_34_elements(193)); -- 
    cr_1513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(193), ack => RPIPE_ConvTranspose_input_pipe_782_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/rr
      -- 
    ca_1514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_782_inst_ack_1, ack => convTranspose_CP_34_elements(194)); -- 
    rr_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => type_cast_786_inst_req_0); -- 
    rr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => RPIPE_ConvTranspose_input_pipe_800_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/ra
      -- 
    ra_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_786_inst_ack_0, ack => convTranspose_CP_34_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	482 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/ca
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_786_inst_ack_1, ack => convTranspose_CP_34_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_update_start_
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/cr
      -- 
    ra_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_800_inst_ack_0, ack => convTranspose_CP_34_elements(197)); -- 
    cr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(197), ack => RPIPE_ConvTranspose_input_pipe_800_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/rr
      -- 
    ca_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_800_inst_ack_1, ack => convTranspose_CP_34_elements(198)); -- 
    rr_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => type_cast_804_inst_req_0); -- 
    rr_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => RPIPE_ConvTranspose_input_pipe_818_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/ra
      -- 
    ra_1551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_0, ack => convTranspose_CP_34_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	482 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/ca
      -- 
    ca_1556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_1, ack => convTranspose_CP_34_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_update_start_
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/cr
      -- 
    ra_1565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_818_inst_ack_0, ack => convTranspose_CP_34_elements(201)); -- 
    cr_1569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(201), ack => RPIPE_ConvTranspose_input_pipe_818_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/rr
      -- 
    ca_1570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_818_inst_ack_1, ack => convTranspose_CP_34_elements(202)); -- 
    rr_1578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(202), ack => type_cast_822_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/ra
      -- 
    ra_1579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_0, ack => convTranspose_CP_34_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	482 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/ca
      -- 
    ca_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_1, ack => convTranspose_CP_34_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/rr
      -- 
    rr_1622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(205), ack => ptr_deref_830_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(172) & convTranspose_CP_34_elements(176) & convTranspose_CP_34_elements(180) & convTranspose_CP_34_elements(184) & convTranspose_CP_34_elements(188) & convTranspose_CP_34_elements(192) & convTranspose_CP_34_elements(196) & convTranspose_CP_34_elements(200) & convTranspose_CP_34_elements(204);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/ra
      -- 
    ra_1623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_830_store_0_ack_0, ack => convTranspose_CP_34_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	482 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_830_store_0_ack_1, ack => convTranspose_CP_34_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	169 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843__exit__
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844__entry__
      -- CP-element group 208: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/$exit
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_38/R_exitcond2_845_place
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_else_link/$entry
      -- 
    branch_req_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(208), ack => if_stmt_844_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(169) & convTranspose_CP_34_elements(207);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	483 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850__exit__
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_38/if_stmt_844_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/if_stmt_844_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_844_branch_ack_1, ack => convTranspose_CP_34_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	478 
    -- CP-element group 210: 	479 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_38/if_stmt_844_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_38/if_stmt_844_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_844_branch_ack_0, ack => convTranspose_CP_34_elements(210)); -- 
    rr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_687_inst_req_0); -- 
    cr_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_687_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	483 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/ra
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_0, ack => convTranspose_CP_34_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	483 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/ca
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_1, ack => convTranspose_CP_34_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	483 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_0, ack => convTranspose_CP_34_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	483 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_1, ack => convTranspose_CP_34_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	483 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => convTranspose_CP_34_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	483 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_1, ack => convTranspose_CP_34_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: 	212 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880__exit__
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881__entry__
      -- CP-element group 217: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/$exit
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_38/R_cmp264505_882_place
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_else_link/$entry
      -- 
    branch_req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(217), ack => if_stmt_881_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(214) & convTranspose_CP_34_elements(216) & convTranspose_CP_34_elements(212);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887__exit__
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922__entry__
      -- CP-element group 218: 	 branch_block_stmt_38/if_stmt_881_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/if_stmt_881_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_update_start_
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/dummy
      -- 
    if_choice_transition_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_881_branch_ack_1, ack => convTranspose_CP_34_elements(218)); -- 
    rr_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_908_inst_req_0); -- 
    cr_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_908_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	490 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_38/if_stmt_881_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_38/if_stmt_881_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_881_branch_ack_0, ack => convTranspose_CP_34_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/ra
      -- 
    ra_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_0, ack => convTranspose_CP_34_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	484 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922__exit__
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/$exit
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/$entry
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$entry
      -- 
    ca_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_1, ack => convTranspose_CP_34_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	489 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/ack
      -- 
    ack_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_937_index_offset_ack_0, ack => convTranspose_CP_34_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	489 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/req
      -- 
    ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_937_index_offset_ack_1, ack => convTranspose_CP_34_elements(223)); -- 
    req_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(223), ack => addr_of_938_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/ack
      -- 
    ack_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_938_final_reg_ack_0, ack => convTranspose_CP_34_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	489 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/rr
      -- 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_938_final_reg_ack_1, ack => convTranspose_CP_34_elements(225)); -- 
    rr_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(225), ack => ptr_deref_941_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/ra
      -- 
    ra_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_0, ack => convTranspose_CP_34_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	489 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/ca
      -- 
    ca_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_1, ack => convTranspose_CP_34_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955__exit__
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956__entry__
      -- CP-element group 228: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_38/R_exitcond_957_place
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_else_link/$entry
      -- 
    branch_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(228), ack => if_stmt_956_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(222) & convTranspose_CP_34_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	490 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962__exit__
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_38/if_stmt_956_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/if_stmt_956_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_1, ack => convTranspose_CP_34_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	485 
    -- CP-element group 230: 	486 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_38/if_stmt_956_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_38/if_stmt_956_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_0, ack => convTranspose_CP_34_elements(230)); -- 
    rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_928_inst_req_0); -- 
    cr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_928_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	490 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/cra
      -- 
    cra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_967_call_ack_0, ack => convTranspose_CP_34_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	490 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/rr
      -- 
    cca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_967_call_ack_1, ack => convTranspose_CP_34_elements(232)); -- 
    rr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(232), ack => type_cast_972_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/ra
      -- 
    ra_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_0, ack => convTranspose_CP_34_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	490 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234: 	349 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234:  members (55) 
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973__exit__
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186__entry__
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/$exit
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/cr
      -- 
    ca_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_1, ack => convTranspose_CP_34_elements(234)); -- 
    req_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    cr_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1054_inst_req_1); -- 
    rr_2216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1054_inst_req_0); -- 
    req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block2_start_1075_inst_req_0); -- 
    cr_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1061_inst_req_1); -- 
    rr_2244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1061_inst_req_0); -- 
    req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block0_start_975_inst_req_0); -- 
    rr_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1110_inst_req_0); -- 
    cr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1110_inst_req_1); -- 
    rr_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1117_inst_req_0); -- 
    cr_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1117_inst_req_1); -- 
    req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block3_start_1131_inst_req_0); -- 
    rr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1166_inst_req_0); -- 
    cr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1166_inst_req_1); -- 
    rr_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1173_inst_req_0); -- 
    cr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1173_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_update_start_
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/req
      -- 
    ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_0, ack => convTranspose_CP_34_elements(235)); -- 
    req_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(235), ack => WPIPE_Block0_start_975_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_975_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_sample_start_
      -- 
    ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_1, ack => convTranspose_CP_34_elements(236)); -- 
    req_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(236), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/req
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_update_start_
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_sample_completed_
      -- 
    ack_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_34_elements(237)); -- 
    req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(237), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_978_update_completed_
      -- 
    ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_34_elements(238)); -- 
    req_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(238), ack => WPIPE_Block0_start_981_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_update_start_
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/req
      -- 
    ack_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_0, ack => convTranspose_CP_34_elements(239)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(239), ack => WPIPE_Block0_start_981_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/req
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_981_Update/$exit
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_1, ack => convTranspose_CP_34_elements(240)); -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(240), ack => WPIPE_Block0_start_984_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/req
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_update_start_
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_sample_completed_
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_0, ack => convTranspose_CP_34_elements(241)); -- 
    req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(241), ack => WPIPE_Block0_start_984_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_984_update_completed_
      -- 
    ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_1, ack => convTranspose_CP_34_elements(242)); -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(242), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_update_start_
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/req
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Sample/$exit
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_34_elements(243)); -- 
    req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(243), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/$entry
      -- 
    ack_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_34_elements(244)); -- 
    req_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(244), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_update_start_
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/req
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Sample/$exit
      -- 
    ack_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_34_elements(245)); -- 
    req_1969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(245), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_990_update_completed_
      -- 
    ack_1970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_34_elements(246)); -- 
    req_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(246), ack => WPIPE_Block0_start_993_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/req
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_update_start_
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_sample_completed_
      -- 
    ack_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_0, ack => convTranspose_CP_34_elements(247)); -- 
    req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(247), ack => WPIPE_Block0_start_993_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_993_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/req
      -- 
    ack_1984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_1, ack => convTranspose_CP_34_elements(248)); -- 
    req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(248), ack => WPIPE_Block0_start_996_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_update_start_
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/req
      -- 
    ack_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_0, ack => convTranspose_CP_34_elements(249)); -- 
    req_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(249), ack => WPIPE_Block0_start_996_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_996_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/req
      -- 
    ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_1, ack => convTranspose_CP_34_elements(250)); -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(250), ack => WPIPE_Block0_start_999_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_update_start_
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/req
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Sample/$exit
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_999_inst_ack_0, ack => convTranspose_CP_34_elements(251)); -- 
    req_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(251), ack => WPIPE_Block0_start_999_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_999_Update/$exit
      -- 
    ack_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_999_inst_ack_1, ack => convTranspose_CP_34_elements(252)); -- 
    req_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(252), ack => WPIPE_Block0_start_1002_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_update_start_
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/req
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_sample_completed_
      -- 
    ack_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_0, ack => convTranspose_CP_34_elements(253)); -- 
    req_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(253), ack => WPIPE_Block0_start_1002_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1002_Update/ack
      -- 
    ack_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_1, ack => convTranspose_CP_34_elements(254)); -- 
    req_2034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(254), ack => WPIPE_Block0_start_1006_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/req
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_update_start_
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_sample_completed_
      -- 
    ack_2035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_0, ack => convTranspose_CP_34_elements(255)); -- 
    req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(255), ack => WPIPE_Block0_start_1006_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1006_update_completed_
      -- 
    ack_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_1, ack => convTranspose_CP_34_elements(256)); -- 
    req_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(256), ack => WPIPE_Block0_start_1010_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/req
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_update_start_
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_sample_completed_
      -- 
    ack_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_0, ack => convTranspose_CP_34_elements(257)); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(257), ack => WPIPE_Block0_start_1010_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1010_update_completed_
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_1, ack => convTranspose_CP_34_elements(258)); -- 
    req_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(258), ack => WPIPE_Block0_start_1013_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/req
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_update_start_
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_sample_completed_
      -- 
    ack_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1013_inst_ack_0, ack => convTranspose_CP_34_elements(259)); -- 
    req_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(259), ack => WPIPE_Block0_start_1013_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1013_update_completed_
      -- 
    ack_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1013_inst_ack_1, ack => convTranspose_CP_34_elements(260)); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(260), ack => WPIPE_Block0_start_1016_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_update_start_
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/req
      -- 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1016_inst_ack_0, ack => convTranspose_CP_34_elements(261)); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(261), ack => WPIPE_Block0_start_1016_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	365 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block0_start_1016_update_completed_
      -- 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1016_inst_ack_1, ack => convTranspose_CP_34_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_update_start_
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/req
      -- 
    ack_2091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_34_elements(263)); -- 
    req_2095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(263), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/req
      -- 
    ack_2096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_34_elements(264)); -- 
    req_2104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/req
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/$entry
      -- 
    ack_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_34_elements(265)); -- 
    req_2109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(265), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1022_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/req
      -- 
    ack_2110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_34_elements(266)); -- 
    req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(266), ack => WPIPE_Block1_start_1025_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_update_start_
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/req
      -- 
    ack_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_0, ack => convTranspose_CP_34_elements(267)); -- 
    req_2123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(267), ack => WPIPE_Block1_start_1025_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1025_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/$entry
      -- 
    ack_2124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_1, ack => convTranspose_CP_34_elements(268)); -- 
    req_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => WPIPE_Block1_start_1028_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/req
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_update_start_
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_sample_completed_
      -- 
    ack_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_0, ack => convTranspose_CP_34_elements(269)); -- 
    req_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(269), ack => WPIPE_Block1_start_1028_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1028_update_completed_
      -- 
    ack_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_1, ack => convTranspose_CP_34_elements(270)); -- 
    req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(270), ack => WPIPE_Block1_start_1031_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/req
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_update_start_
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_sample_completed_
      -- 
    ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_0, ack => convTranspose_CP_34_elements(271)); -- 
    req_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(271), ack => WPIPE_Block1_start_1031_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1031_update_completed_
      -- 
    ack_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_1, ack => convTranspose_CP_34_elements(272)); -- 
    req_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(272), ack => WPIPE_Block1_start_1034_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/req
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_update_start_
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Sample/ack
      -- 
    ack_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_0, ack => convTranspose_CP_34_elements(273)); -- 
    req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(273), ack => WPIPE_Block1_start_1034_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1034_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/$entry
      -- 
    ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_1, ack => convTranspose_CP_34_elements(274)); -- 
    req_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(274), ack => WPIPE_Block1_start_1037_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_update_start_
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/req
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Sample/$exit
      -- 
    ack_2175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_0, ack => convTranspose_CP_34_elements(275)); -- 
    req_2179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(275), ack => WPIPE_Block1_start_1037_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1037_Update/$exit
      -- 
    ack_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_1, ack => convTranspose_CP_34_elements(276)); -- 
    req_2188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(276), ack => WPIPE_Block1_start_1040_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/req
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_update_start_
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_sample_completed_
      -- 
    ack_2189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1040_inst_ack_0, ack => convTranspose_CP_34_elements(277)); -- 
    req_2193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(277), ack => WPIPE_Block1_start_1040_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1040_update_completed_
      -- 
    ack_2194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1040_inst_ack_1, ack => convTranspose_CP_34_elements(278)); -- 
    req_2202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(278), ack => WPIPE_Block1_start_1043_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/req
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_update_start_
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_sample_completed_
      -- 
    ack_2203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1043_inst_ack_0, ack => convTranspose_CP_34_elements(279)); -- 
    req_2207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(279), ack => WPIPE_Block1_start_1043_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1043_update_completed_
      -- 
    ack_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1043_inst_ack_1, ack => convTranspose_CP_34_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_sample_completed_
      -- 
    ra_2217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_0, ack => convTranspose_CP_34_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1054_update_completed_
      -- 
    ca_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_1, ack => convTranspose_CP_34_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_sample_start_
      -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(283), ack => WPIPE_Block1_start_1056_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(280) & convTranspose_CP_34_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_update_start_
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/req
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_sample_completed_
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_0, ack => convTranspose_CP_34_elements(284)); -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(284), ack => WPIPE_Block1_start_1056_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1056_Update/ack
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_1, ack => convTranspose_CP_34_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_sample_completed_
      -- 
    ra_2245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_0, ack => convTranspose_CP_34_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1061_update_completed_
      -- 
    ca_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_1, ack => convTranspose_CP_34_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_sample_start_
      -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(288), ack => WPIPE_Block1_start_1063_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(285) & convTranspose_CP_34_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_update_start_
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/req
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_sample_completed_
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_0, ack => convTranspose_CP_34_elements(289)); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(289), ack => WPIPE_Block1_start_1063_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1063_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_sample_start_
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_1, ack => convTranspose_CP_34_elements(290)); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(290), ack => WPIPE_Block1_start_1066_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/req
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_update_start_
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_sample_completed_
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_0, ack => convTranspose_CP_34_elements(291)); -- 
    req_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(291), ack => WPIPE_Block1_start_1066_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1066_update_completed_
      -- 
    ack_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_1, ack => convTranspose_CP_34_elements(292)); -- 
    req_2286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(292), ack => WPIPE_Block1_start_1069_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_update_start_
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/req
      -- 
    ack_2287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1069_inst_ack_0, ack => convTranspose_CP_34_elements(293)); -- 
    req_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(293), ack => WPIPE_Block1_start_1069_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1069_Update/ack
      -- 
    ack_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1069_inst_ack_1, ack => convTranspose_CP_34_elements(294)); -- 
    req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(294), ack => WPIPE_Block1_start_1072_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/req
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_update_start_
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_sample_completed_
      -- 
    ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1072_inst_ack_0, ack => convTranspose_CP_34_elements(295)); -- 
    req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(295), ack => WPIPE_Block1_start_1072_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	365 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block1_start_1072_update_completed_
      -- 
    ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1072_inst_ack_1, ack => convTranspose_CP_34_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/req
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_update_start_
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_sample_completed_
      -- 
    ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_0, ack => convTranspose_CP_34_elements(297)); -- 
    req_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(297), ack => WPIPE_Block2_start_1075_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1075_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_sample_start_
      -- 
    ack_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_1, ack => convTranspose_CP_34_elements(298)); -- 
    req_2328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(298), ack => WPIPE_Block2_start_1078_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/req
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_update_start_
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_sample_completed_
      -- 
    ack_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_0, ack => convTranspose_CP_34_elements(299)); -- 
    req_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(299), ack => WPIPE_Block2_start_1078_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1078_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_sample_start_
      -- 
    ack_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_1, ack => convTranspose_CP_34_elements(300)); -- 
    req_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(300), ack => WPIPE_Block2_start_1081_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/req
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_update_start_
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_sample_completed_
      -- 
    ack_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_0, ack => convTranspose_CP_34_elements(301)); -- 
    req_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(301), ack => WPIPE_Block2_start_1081_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1081_update_completed_
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_1, ack => convTranspose_CP_34_elements(302)); -- 
    req_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(302), ack => WPIPE_Block2_start_1084_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/req
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_update_start_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_sample_completed_
      -- 
    ack_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_0, ack => convTranspose_CP_34_elements(303)); -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(303), ack => WPIPE_Block2_start_1084_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1084_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/$entry
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_1, ack => convTranspose_CP_34_elements(304)); -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(304), ack => WPIPE_Block2_start_1087_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_update_start_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/req
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Sample/$exit
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_0, ack => convTranspose_CP_34_elements(305)); -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(305), ack => WPIPE_Block2_start_1087_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1087_update_completed_
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_1, ack => convTranspose_CP_34_elements(306)); -- 
    req_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(306), ack => WPIPE_Block2_start_1090_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_update_start_
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/req
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/$entry
      -- 
    ack_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_0, ack => convTranspose_CP_34_elements(307)); -- 
    req_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(307), ack => WPIPE_Block2_start_1090_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1090_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/req
      -- 
    ack_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_1, ack => convTranspose_CP_34_elements(308)); -- 
    req_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(308), ack => WPIPE_Block2_start_1093_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_update_start_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/req
      -- 
    ack_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_0, ack => convTranspose_CP_34_elements(309)); -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(309), ack => WPIPE_Block2_start_1093_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1093_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/req
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_1, ack => convTranspose_CP_34_elements(310)); -- 
    req_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(310), ack => WPIPE_Block2_start_1096_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_update_start_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/req
      -- 
    ack_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1096_inst_ack_0, ack => convTranspose_CP_34_elements(311)); -- 
    req_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(311), ack => WPIPE_Block2_start_1096_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1096_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/req
      -- 
    ack_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1096_inst_ack_1, ack => convTranspose_CP_34_elements(312)); -- 
    req_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(312), ack => WPIPE_Block2_start_1099_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_update_start_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/req
      -- 
    ack_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1099_inst_ack_0, ack => convTranspose_CP_34_elements(313)); -- 
    req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(313), ack => WPIPE_Block2_start_1099_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1099_Update/ack
      -- 
    ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1099_inst_ack_1, ack => convTranspose_CP_34_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Sample/ra
      -- 
    ra_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => convTranspose_CP_34_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1110_Update/ca
      -- 
    ca_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => convTranspose_CP_34_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/req
      -- 
    req_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => WPIPE_Block2_start_1112_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(314) & convTranspose_CP_34_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_update_start_
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/req
      -- 
    ack_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1112_inst_ack_0, ack => convTranspose_CP_34_elements(318)); -- 
    req_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(318), ack => WPIPE_Block2_start_1112_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1112_Update/ack
      -- 
    ack_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1112_inst_ack_1, ack => convTranspose_CP_34_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Sample/ra
      -- 
    ra_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1117_inst_ack_0, ack => convTranspose_CP_34_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1117_Update/ca
      -- 
    ca_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1117_inst_ack_1, ack => convTranspose_CP_34_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/req
      -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(322), ack => WPIPE_Block2_start_1119_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(319) & convTranspose_CP_34_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_update_start_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/req
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_0, ack => convTranspose_CP_34_elements(323)); -- 
    req_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(323), ack => WPIPE_Block2_start_1119_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1119_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/req
      -- 
    ack_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_1, ack => convTranspose_CP_34_elements(324)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(324), ack => WPIPE_Block2_start_1122_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_update_start_
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/req
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_0, ack => convTranspose_CP_34_elements(325)); -- 
    req_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(325), ack => WPIPE_Block2_start_1122_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1122_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/req
      -- 
    ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_1, ack => convTranspose_CP_34_elements(326)); -- 
    req_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(326), ack => WPIPE_Block2_start_1125_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_update_start_
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/req
      -- 
    ack_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_0, ack => convTranspose_CP_34_elements(327)); -- 
    req_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(327), ack => WPIPE_Block2_start_1125_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1125_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/req
      -- 
    ack_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_1, ack => convTranspose_CP_34_elements(328)); -- 
    req_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(328), ack => WPIPE_Block2_start_1128_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_update_start_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/req
      -- 
    ack_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_0, ack => convTranspose_CP_34_elements(329)); -- 
    req_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(329), ack => WPIPE_Block2_start_1128_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	365 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block2_start_1128_Update/ack
      -- 
    ack_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_1, ack => convTranspose_CP_34_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_update_start_
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/req
      -- 
    ack_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_0, ack => convTranspose_CP_34_elements(331)); -- 
    req_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(331), ack => WPIPE_Block3_start_1131_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1131_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/req
      -- 
    ack_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_1, ack => convTranspose_CP_34_elements(332)); -- 
    req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(332), ack => WPIPE_Block3_start_1134_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_update_start_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/req
      -- 
    ack_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_0, ack => convTranspose_CP_34_elements(333)); -- 
    req_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(333), ack => WPIPE_Block3_start_1134_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1134_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/req
      -- 
    ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_1, ack => convTranspose_CP_34_elements(334)); -- 
    req_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(334), ack => WPIPE_Block3_start_1137_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_update_start_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/req
      -- 
    ack_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_0, ack => convTranspose_CP_34_elements(335)); -- 
    req_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(335), ack => WPIPE_Block3_start_1137_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1137_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/req
      -- 
    ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_1, ack => convTranspose_CP_34_elements(336)); -- 
    req_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(336), ack => WPIPE_Block3_start_1140_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_update_start_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/req
      -- 
    ack_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_0, ack => convTranspose_CP_34_elements(337)); -- 
    req_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(337), ack => WPIPE_Block3_start_1140_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1140_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/req
      -- 
    ack_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_1, ack => convTranspose_CP_34_elements(338)); -- 
    req_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(338), ack => WPIPE_Block3_start_1143_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_update_start_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/req
      -- 
    ack_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_0, ack => convTranspose_CP_34_elements(339)); -- 
    req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(339), ack => WPIPE_Block3_start_1143_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1143_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/req
      -- 
    ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_1, ack => convTranspose_CP_34_elements(340)); -- 
    req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(340), ack => WPIPE_Block3_start_1146_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_update_start_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/req
      -- 
    ack_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_0, ack => convTranspose_CP_34_elements(341)); -- 
    req_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(341), ack => WPIPE_Block3_start_1146_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1146_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/req
      -- 
    ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_1, ack => convTranspose_CP_34_elements(342)); -- 
    req_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(342), ack => WPIPE_Block3_start_1149_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_update_start_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/req
      -- 
    ack_2623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_0, ack => convTranspose_CP_34_elements(343)); -- 
    req_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(343), ack => WPIPE_Block3_start_1149_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1149_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/req
      -- 
    ack_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_1, ack => convTranspose_CP_34_elements(344)); -- 
    req_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(344), ack => WPIPE_Block3_start_1152_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_update_start_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/req
      -- 
    ack_2637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1152_inst_ack_0, ack => convTranspose_CP_34_elements(345)); -- 
    req_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(345), ack => WPIPE_Block3_start_1152_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1152_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/req
      -- 
    ack_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1152_inst_ack_1, ack => convTranspose_CP_34_elements(346)); -- 
    req_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(346), ack => WPIPE_Block3_start_1155_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_update_start_
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/req
      -- 
    ack_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1155_inst_ack_0, ack => convTranspose_CP_34_elements(347)); -- 
    req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(347), ack => WPIPE_Block3_start_1155_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1155_Update/ack
      -- 
    ack_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1155_inst_ack_1, ack => convTranspose_CP_34_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Sample/ra
      -- 
    ra_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_0, ack => convTranspose_CP_34_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1166_Update/ca
      -- 
    ca_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_1, ack => convTranspose_CP_34_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/req
      -- 
    req_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(351), ack => WPIPE_Block3_start_1168_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(348) & convTranspose_CP_34_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_update_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/req
      -- 
    ack_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1168_inst_ack_0, ack => convTranspose_CP_34_elements(352)); -- 
    req_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(352), ack => WPIPE_Block3_start_1168_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1168_Update/ack
      -- 
    ack_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1168_inst_ack_1, ack => convTranspose_CP_34_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Sample/ra
      -- 
    ra_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => convTranspose_CP_34_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/type_cast_1173_Update/ca
      -- 
    ca_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => convTranspose_CP_34_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/req
      -- 
    req_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(356), ack => WPIPE_Block3_start_1175_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(353) & convTranspose_CP_34_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_update_start_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/req
      -- 
    ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_0, ack => convTranspose_CP_34_elements(357)); -- 
    req_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(357), ack => WPIPE_Block3_start_1175_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1175_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/req
      -- 
    ack_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_1, ack => convTranspose_CP_34_elements(358)); -- 
    req_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(358), ack => WPIPE_Block3_start_1178_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_update_start_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/req
      -- 
    ack_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_0, ack => convTranspose_CP_34_elements(359)); -- 
    req_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(359), ack => WPIPE_Block3_start_1178_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1178_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/req
      -- 
    ack_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_1, ack => convTranspose_CP_34_elements(360)); -- 
    req_2734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(360), ack => WPIPE_Block3_start_1181_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_update_start_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/req
      -- 
    ack_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_0, ack => convTranspose_CP_34_elements(361)); -- 
    req_2739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(361), ack => WPIPE_Block3_start_1181_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1181_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/req
      -- 
    ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_1, ack => convTranspose_CP_34_elements(362)); -- 
    req_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(362), ack => WPIPE_Block3_start_1184_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_update_start_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/req
      -- 
    ack_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_0, ack => convTranspose_CP_34_elements(363)); -- 
    req_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(363), ack => WPIPE_Block3_start_1184_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/WPIPE_Block3_start_1184_Update/ack
      -- 
    ack_2754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_1, ack => convTranspose_CP_34_elements(364)); -- 
    -- CP-element group 365:  join  fork  transition  place  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	262 
    -- CP-element group 365: 	296 
    -- CP-element group 365: 	364 
    -- CP-element group 365: 	330 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: 	368 
    -- CP-element group 365: 	370 
    -- CP-element group 365: 	372 
    -- CP-element group 365:  members (16) 
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186__exit__
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199__entry__
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1186/$exit
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/rr
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/rr
      -- 
    rr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block0_done_1189_inst_req_0); -- 
    rr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block1_done_1192_inst_req_0); -- 
    rr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block2_done_1195_inst_req_0); -- 
    rr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block3_done_1198_inst_req_0); -- 
    convTranspose_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(262) & convTranspose_CP_34_elements(296) & convTranspose_CP_34_elements(364) & convTranspose_CP_34_elements(330);
      gj_convTranspose_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (6) 
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_update_start_
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Sample/ra
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/cr
      -- 
    ra_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1189_inst_ack_0, ack => convTranspose_CP_34_elements(366)); -- 
    cr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(366), ack => RPIPE_Block0_done_1189_inst_req_1); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	374 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block0_done_1189_Update/ca
      -- 
    ca_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1189_inst_ack_1, ack => convTranspose_CP_34_elements(367)); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	365 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_update_start_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Sample/ra
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/cr
      -- 
    ra_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1192_inst_ack_0, ack => convTranspose_CP_34_elements(368)); -- 
    cr_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(368), ack => RPIPE_Block1_done_1192_inst_req_1); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block1_done_1192_Update/ca
      -- 
    ca_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1192_inst_ack_1, ack => convTranspose_CP_34_elements(369)); -- 
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_update_start_
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Sample/ra
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/cr
      -- 
    ra_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1195_inst_ack_0, ack => convTranspose_CP_34_elements(370)); -- 
    cr_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(370), ack => RPIPE_Block2_done_1195_inst_req_1); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	374 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block2_done_1195_Update/ca
      -- 
    ca_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1195_inst_ack_1, ack => convTranspose_CP_34_elements(371)); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	365 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_update_start_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Sample/ra
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/cr
      -- 
    ra_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1198_inst_ack_0, ack => convTranspose_CP_34_elements(372)); -- 
    cr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(372), ack => RPIPE_Block3_done_1198_inst_req_1); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/RPIPE_Block3_done_1198_Update/ca
      -- 
    ca_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1198_inst_ack_1, ack => convTranspose_CP_34_elements(373)); -- 
    -- CP-element group 374:  join  fork  transition  place  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	367 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	371 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	388 
    -- CP-element group 374: 	390 
    -- CP-element group 374: 	392 
    -- CP-element group 374: 	394 
    -- CP-element group 374: 	384 
    -- CP-element group 374: 	386 
    -- CP-element group 374: 	375 
    -- CP-element group 374: 	376 
    -- CP-element group 374: 	378 
    -- CP-element group 374: 	380 
    -- CP-element group 374: 	382 
    -- CP-element group 374:  members (37) 
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199__exit__
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310__entry__
      -- CP-element group 374: 	 branch_block_stmt_38/assign_stmt_1190_to_assign_stmt_1199/$exit
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/crr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/ccr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_update_start_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/cr
      -- 
    crr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => call_stmt_1202_call_req_0); -- 
    ccr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => call_stmt_1202_call_req_1); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1206_inst_req_1); -- 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1215_inst_req_1); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1225_inst_req_1); -- 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1235_inst_req_1); -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1245_inst_req_1); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1255_inst_req_1); -- 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1265_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1275_inst_req_1); -- 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(374), ack => type_cast_1285_inst_req_1); -- 
    convTranspose_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(367) & convTranspose_CP_34_elements(369) & convTranspose_CP_34_elements(371) & convTranspose_CP_34_elements(373);
      gj_convTranspose_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Sample/cra
      -- 
    cra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1202_call_ack_0, ack => convTranspose_CP_34_elements(375)); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/call_stmt_1202_Update/cca
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/rr
      -- 
    cca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1202_call_ack_1, ack => convTranspose_CP_34_elements(376)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(376), ack => type_cast_1206_inst_req_0); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_0, ack => convTranspose_CP_34_elements(377)); -- 
    -- CP-element group 378:  fork  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	374 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	387 
    -- CP-element group 378: 	389 
    -- CP-element group 378: 	391 
    -- CP-element group 378: 	393 
    -- CP-element group 378: 	383 
    -- CP-element group 378: 	385 
    -- CP-element group 378: 	379 
    -- CP-element group 378: 	381 
    -- CP-element group 378:  members (27) 
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1206_Update/ca
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/rr
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/rr
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1206_inst_ack_1, ack => convTranspose_CP_34_elements(378)); -- 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1265_inst_req_0); -- 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1275_inst_req_0); -- 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1285_inst_req_0); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1235_inst_req_0); -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1245_inst_req_0); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1255_inst_req_0); -- 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1215_inst_req_0); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(378), ack => type_cast_1225_inst_req_0); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Sample/ra
      -- 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_0, ack => convTranspose_CP_34_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	374 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	415 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1215_Update/ca
      -- 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_1, ack => convTranspose_CP_34_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	378 
    -- CP-element group 381: successors 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Sample/ra
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1225_inst_ack_0, ack => convTranspose_CP_34_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	374 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	412 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1225_Update/ca
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1225_inst_ack_1, ack => convTranspose_CP_34_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	378 
    -- CP-element group 383: successors 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_sample_completed_
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Sample/ra
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_0, ack => convTranspose_CP_34_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	374 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	409 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_update_completed_
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1235_Update/ca
      -- 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1235_inst_ack_1, ack => convTranspose_CP_34_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	378 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Sample/ra
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1245_inst_ack_0, ack => convTranspose_CP_34_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	374 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	406 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1245_Update/ca
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1245_inst_ack_1, ack => convTranspose_CP_34_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	378 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_0, ack => convTranspose_CP_34_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	374 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	403 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1255_Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_1, ack => convTranspose_CP_34_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	378 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Sample/ra
      -- 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_0, ack => convTranspose_CP_34_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	374 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	400 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1265_Update/ca
      -- 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_1, ack => convTranspose_CP_34_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	378 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Sample/ra
      -- 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_0, ack => convTranspose_CP_34_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	374 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	397 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1275_Update/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1275_inst_ack_1, ack => convTranspose_CP_34_elements(392)); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	378 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/$exit
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Sample/ra
      -- 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1285_inst_ack_0, ack => convTranspose_CP_34_elements(393)); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	374 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/$exit
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/type_cast_1285_Update/ca
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_sample_start_
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/req
      -- 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1285_inst_ack_1, ack => convTranspose_CP_34_elements(394)); -- 
    req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(394), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_0); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/req
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_update_start_
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Sample/ack
      -- 
    ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0, ack => convTranspose_CP_34_elements(395)); -- 
    req_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(395), ack => WPIPE_ConvTranspose_output_pipe_1287_inst_req_1); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_Update/ack
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1287_update_completed_
      -- 
    ack_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1, ack => convTranspose_CP_34_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	392 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/req
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/$entry
      -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(397), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_0); -- 
    convTranspose_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(392) & convTranspose_CP_34_elements(396);
      gj_convTranspose_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  transition  input  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (6) 
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Sample/ack
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_update_start_
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/req
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0, ack => convTranspose_CP_34_elements(398)); -- 
    req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(398), ack => WPIPE_ConvTranspose_output_pipe_1290_inst_req_1); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1290_Update/ack
      -- 
    ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1, ack => convTranspose_CP_34_elements(399)); -- 
    -- CP-element group 400:  join  transition  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	390 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/req
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_sample_start_
      -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(400), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_0); -- 
    convTranspose_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(390) & convTranspose_CP_34_elements(399);
      gj_convTranspose_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  transition  input  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (6) 
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/req
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/ack
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_update_start_
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_sample_completed_
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0, ack => convTranspose_CP_34_elements(401)); -- 
    req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(401), ack => WPIPE_ConvTranspose_output_pipe_1293_inst_req_1); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/ack
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1293_update_completed_
      -- 
    ack_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1, ack => convTranspose_CP_34_elements(402)); -- 
    -- CP-element group 403:  join  transition  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	388 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/req
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_sample_start_
      -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_0); -- 
    convTranspose_cp_element_group_403: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_403"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(388) & convTranspose_CP_34_elements(402);
      gj_convTranspose_cp_element_group_403 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(403), clk => clk, reset => reset); --
    end block;
    -- CP-element group 404:  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (6) 
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/req
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/ack
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_update_start_
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_sample_completed_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0, ack => convTranspose_CP_34_elements(404)); -- 
    req_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(404), ack => WPIPE_ConvTranspose_output_pipe_1296_inst_req_1); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/ack
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1296_update_completed_
      -- 
    ack_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1, ack => convTranspose_CP_34_elements(405)); -- 
    -- CP-element group 406:  join  transition  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: 	386 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/req
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_sample_start_
      -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_0); -- 
    convTranspose_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(405) & convTranspose_CP_34_elements(386);
      gj_convTranspose_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  transition  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (6) 
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/req
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Sample/ack
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_update_start_
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_sample_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0, ack => convTranspose_CP_34_elements(407)); -- 
    req_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(407), ack => WPIPE_ConvTranspose_output_pipe_1299_inst_req_1); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/ack
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1299_update_completed_
      -- 
    ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1, ack => convTranspose_CP_34_elements(408)); -- 
    -- CP-element group 409:  join  transition  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: 	384 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/req
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/$entry
      -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_0); -- 
    convTranspose_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(408) & convTranspose_CP_34_elements(384);
      gj_convTranspose_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (6) 
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/req
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_update_start_
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Sample/ack
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0, ack => convTranspose_CP_34_elements(410)); -- 
    req_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(410), ack => WPIPE_ConvTranspose_output_pipe_1302_inst_req_1); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1302_Update/ack
      -- 
    ack_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1, ack => convTranspose_CP_34_elements(411)); -- 
    -- CP-element group 412:  join  transition  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: 	382 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/$entry
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_sample_start_
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/req
      -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1305_inst_req_0); -- 
    convTranspose_cp_element_group_412: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_412"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(411) & convTranspose_CP_34_elements(382);
      gj_convTranspose_cp_element_group_412 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(412), clk => clk, reset => reset); --
    end block;
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (6) 
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_update_start_
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_sample_completed_
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/req
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/$entry
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/ack
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Sample/$exit
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1305_inst_ack_0, ack => convTranspose_CP_34_elements(413)); -- 
    req_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(413), ack => WPIPE_ConvTranspose_output_pipe_1305_inst_req_1); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_update_completed_
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/ack
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1305_Update/$exit
      -- 
    ack_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1305_inst_ack_1, ack => convTranspose_CP_34_elements(414)); -- 
    -- CP-element group 415:  join  transition  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: 	380 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/req
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_sample_start_
      -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1308_inst_req_0); -- 
    convTranspose_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(414) & convTranspose_CP_34_elements(380);
      gj_convTranspose_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/req
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/$entry
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_update_start_
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_sample_completed_
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1308_inst_ack_0, ack => convTranspose_CP_34_elements(416)); -- 
    req_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(416), ack => WPIPE_ConvTranspose_output_pipe_1308_inst_req_1); -- 
    -- CP-element group 417:  branch  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417: 	419 
    -- CP-element group 417:  members (13) 
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310__exit__
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312__entry__
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_else_link/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_if_link/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_eval_test/branch_req
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_eval_test/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_eval_test/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1312_dead_link/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/WPIPE_ConvTranspose_output_pipe_1308_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_38/R_cmp264505_1313_place
      -- CP-element group 417: 	 branch_block_stmt_38/call_stmt_1202_to_assign_stmt_1310/$exit
      -- 
    ack_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1308_inst_ack_1, ack => convTranspose_CP_34_elements(417)); -- 
    branch_req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(417), ack => if_stmt_1312_branch_req_0); -- 
    -- CP-element group 418:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: 	421 
    -- CP-element group 418:  members (18) 
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318__exit__
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353__entry__
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/cr
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/rr
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_update_start_
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/if_stmt_1312_if_link/if_choice_transition
      -- CP-element group 418: 	 branch_block_stmt_38/if_stmt_1312_if_link/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_bbx_xnph
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiReqMerge
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiAck/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiAck/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/merge_stmt_1318_PhiAck/dummy
      -- 
    if_choice_transition_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1312_branch_ack_1, ack => convTranspose_CP_34_elements(418)); -- 
    cr_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(418), ack => type_cast_1339_inst_req_1); -- 
    rr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(418), ack => type_cast_1339_inst_req_0); -- 
    -- CP-element group 419:  transition  place  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	497 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_38/forx_xend273_forx_xend500
      -- CP-element group 419: 	 branch_block_stmt_38/if_stmt_1312_else_link/else_choice_transition
      -- CP-element group 419: 	 branch_block_stmt_38/if_stmt_1312_else_link/$exit
      -- CP-element group 419: 	 branch_block_stmt_38/forx_xend273_forx_xend500_PhiReq/$entry
      -- CP-element group 419: 	 branch_block_stmt_38/forx_xend273_forx_xend500_PhiReq/$exit
      -- 
    else_choice_transition_3085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1312_branch_ack_0, ack => convTranspose_CP_34_elements(419)); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/ra
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_sample_completed_
      -- 
    ra_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_0, ack => convTranspose_CP_34_elements(420)); -- 
    -- CP-element group 421:  transition  place  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	418 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	491 
    -- CP-element group 421:  members (9) 
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353__exit__
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/ca
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/type_cast_1339_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1324_to_assign_stmt_1353/$exit
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/$entry
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/$entry
      -- CP-element group 421: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$entry
      -- 
    ca_3104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1339_inst_ack_1, ack => convTranspose_CP_34_elements(421)); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	496 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	467 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_sample_complete
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/ack
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/$exit
      -- 
    ack_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1368_index_offset_ack_0, ack => convTranspose_CP_34_elements(422)); -- 
    -- CP-element group 423:  transition  input  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	496 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (11) 
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_sample_start_
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_root_address_calculated
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_offset_calculated
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/req
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/$entry
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/sum_rename_ack
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/sum_rename_req
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/$exit
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_base_plus_offset/$entry
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/ack
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/$exit
      -- 
    ack_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1368_index_offset_ack_1, ack => convTranspose_CP_34_elements(423)); -- 
    req_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(423), ack => addr_of_1369_final_reg_req_0); -- 
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/ack
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_request/$exit
      -- 
    ack_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1369_final_reg_ack_0, ack => convTranspose_CP_34_elements(424)); -- 
    -- CP-element group 425:  join  fork  transition  input  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	496 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (24) 
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/rr
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/root_register_ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/root_register_req
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_addrgen/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/sum_rename_ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/sum_rename_req
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_plus_offset/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/base_resize_ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/base_resize_req
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_addr_resize/$entry
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_address_resized
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_root_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_word_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_base_address_calculated
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_sample_start_
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/ack
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/$exit
      -- 
    ack_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1369_final_reg_ack_1, ack => convTranspose_CP_34_elements(425)); -- 
    rr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(425), ack => ptr_deref_1373_load_0_req_0); -- 
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426:  members (5) 
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/ra
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/word_0/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/word_access_start/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_sample_completed_
      -- 
    ra_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1373_load_0_ack_0, ack => convTranspose_CP_34_elements(426)); -- 
    -- CP-element group 427:  fork  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	496 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427: 	430 
    -- CP-element group 427: 	432 
    -- CP-element group 427: 	434 
    -- CP-element group 427: 	436 
    -- CP-element group 427: 	438 
    -- CP-element group 427: 	440 
    -- CP-element group 427: 	442 
    -- CP-element group 427:  members (33) 
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/ca
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/merge_ack
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/merge_req
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/ptr_deref_1373_Merge/$exit
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_sample_start_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/rr
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/$entry
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_sample_start_
      -- 
    ca_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1373_load_0_ack_1, ack => convTranspose_CP_34_elements(427)); -- 
    rr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1377_inst_req_0); -- 
    rr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1387_inst_req_0); -- 
    rr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1397_inst_req_0); -- 
    rr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1407_inst_req_0); -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1417_inst_req_0); -- 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1427_inst_req_0); -- 
    rr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1437_inst_req_0); -- 
    rr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(427), ack => type_cast_1447_inst_req_0); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/ra
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_sample_completed_
      -- 
    ra_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1377_inst_ack_0, ack => convTranspose_CP_34_elements(428)); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	496 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	464 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/ca
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_update_completed_
      -- 
    ca_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1377_inst_ack_1, ack => convTranspose_CP_34_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	427 
    -- CP-element group 430: successors 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/ra
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Sample/$exit
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_sample_completed_
      -- 
    ra_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_0, ack => convTranspose_CP_34_elements(430)); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	496 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	461 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/ca
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/$exit
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_update_completed_
      -- 
    ca_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_1, ack => convTranspose_CP_34_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	427 
    -- CP-element group 432: successors 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Sample/ra
      -- 
    ra_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1397_inst_ack_0, ack => convTranspose_CP_34_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	496 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	458 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/ca
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/$exit
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1397_inst_ack_1, ack => convTranspose_CP_34_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	427 
    -- CP-element group 434: successors 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/ra
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Sample/$exit
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_sample_completed_
      -- 
    ra_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1407_inst_ack_0, ack => convTranspose_CP_34_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	496 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	455 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/ca
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/$exit
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_update_completed_
      -- 
    ca_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1407_inst_ack_1, ack => convTranspose_CP_34_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	427 
    -- CP-element group 436: successors 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/$exit
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Sample/ra
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_sample_completed_
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_0, ack => convTranspose_CP_34_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	496 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	452 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/ca
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_update_completed_
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/$exit
      -- 
    ca_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_1, ack => convTranspose_CP_34_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	427 
    -- CP-element group 438: successors 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/ra
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_sample_completed_
      -- 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_0, ack => convTranspose_CP_34_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	496 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	449 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/ca
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_update_completed_
      -- 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_1, ack => convTranspose_CP_34_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	427 
    -- CP-element group 440: successors 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_sample_completed_
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/ra
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Sample/$exit
      -- 
    ra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_0, ack => convTranspose_CP_34_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	496 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	446 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/ca
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_update_completed_
      -- 
    ca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_1, ack => convTranspose_CP_34_elements(441)); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	427 
    -- CP-element group 442: successors 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/ra
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Sample/$exit
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_sample_completed_
      -- 
    ra_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1447_inst_ack_0, ack => convTranspose_CP_34_elements(442)); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	496 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/req
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/ca
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/$exit
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_update_completed_
      -- 
    ca_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1447_inst_ack_1, ack => convTranspose_CP_34_elements(443)); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(443), ack => WPIPE_ConvTranspose_output_pipe_1449_inst_req_0); -- 
    -- CP-element group 444:  transition  input  output  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (6) 
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/req
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/ack
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_update_start_
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_sample_completed_
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0, ack => convTranspose_CP_34_elements(444)); -- 
    req_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(444), ack => WPIPE_ConvTranspose_output_pipe_1449_inst_req_1); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/ack
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1449_update_completed_
      -- 
    ack_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1, ack => convTranspose_CP_34_elements(445)); -- 
    -- CP-element group 446:  join  transition  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	441 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/req
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_sample_start_
      -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1452_inst_req_0); -- 
    convTranspose_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(441) & convTranspose_CP_34_elements(445);
      gj_convTranspose_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  transition  input  output  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (6) 
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/req
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/$entry
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/ack
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_update_start_
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_sample_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0, ack => convTranspose_CP_34_elements(447)); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(447), ack => WPIPE_ConvTranspose_output_pipe_1452_inst_req_1); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/ack
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1452_update_completed_
      -- 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1, ack => convTranspose_CP_34_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	439 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/req
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/$entry
      -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1455_inst_req_0); -- 
    convTranspose_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(439) & convTranspose_CP_34_elements(448);
      gj_convTranspose_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (6) 
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_update_start_
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/req
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_sample_completed_
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/ack
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Sample/$exit
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0, ack => convTranspose_CP_34_elements(450)); -- 
    req_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(450), ack => WPIPE_ConvTranspose_output_pipe_1455_inst_req_1); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/ack
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1455_update_completed_
      -- 
    ack_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1, ack => convTranspose_CP_34_elements(451)); -- 
    -- CP-element group 452:  join  transition  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	437 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/req
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_sample_start_
      -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1458_inst_req_0); -- 
    convTranspose_cp_element_group_452: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_452"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(437) & convTranspose_CP_34_elements(451);
      gj_convTranspose_cp_element_group_452 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(452), clk => clk, reset => reset); --
    end block;
    -- CP-element group 453:  transition  input  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (6) 
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/req
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/ack
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Sample/$exit
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_update_start_
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_sample_completed_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0, ack => convTranspose_CP_34_elements(453)); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(453), ack => WPIPE_ConvTranspose_output_pipe_1458_inst_req_1); -- 
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/ack
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_Update/$exit
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1458_update_completed_
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1, ack => convTranspose_CP_34_elements(454)); -- 
    -- CP-element group 455:  join  transition  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	435 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_sample_start_
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/req
      -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1461_inst_req_0); -- 
    convTranspose_cp_element_group_455: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_455"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(435) & convTranspose_CP_34_elements(454);
      gj_convTranspose_cp_element_group_455 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 456:  transition  input  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (6) 
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_update_start_
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_sample_completed_
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/$exit
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Sample/ack
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/req
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0, ack => convTranspose_CP_34_elements(456)); -- 
    req_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(456), ack => WPIPE_ConvTranspose_output_pipe_1461_inst_req_1); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_update_completed_
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/$exit
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1461_Update/ack
      -- 
    ack_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1, ack => convTranspose_CP_34_elements(457)); -- 
    -- CP-element group 458:  join  transition  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	433 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_sample_start_
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/req
      -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1464_inst_req_0); -- 
    convTranspose_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(433) & convTranspose_CP_34_elements(457);
      gj_convTranspose_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  transition  input  output  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (6) 
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_update_start_
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Sample/ack
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/$entry
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/req
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0, ack => convTranspose_CP_34_elements(459)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(459), ack => WPIPE_ConvTranspose_output_pipe_1464_inst_req_1); -- 
    -- CP-element group 460:  transition  input  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1464_Update/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1, ack => convTranspose_CP_34_elements(460)); -- 
    -- CP-element group 461:  join  transition  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	431 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/req
      -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1467_inst_req_0); -- 
    convTranspose_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(431) & convTranspose_CP_34_elements(460);
      gj_convTranspose_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  transition  input  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (6) 
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_sample_completed_
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_update_start_
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/$exit
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Sample/ack
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/req
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1467_inst_ack_0, ack => convTranspose_CP_34_elements(462)); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(462), ack => WPIPE_ConvTranspose_output_pipe_1467_inst_req_1); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_update_completed_
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/$exit
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1467_Update/ack
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1467_inst_ack_1, ack => convTranspose_CP_34_elements(463)); -- 
    -- CP-element group 464:  join  transition  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	429 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_sample_start_
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/$entry
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/req
      -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1470_inst_req_0); -- 
    convTranspose_cp_element_group_464: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_464"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(429) & convTranspose_CP_34_elements(463);
      gj_convTranspose_cp_element_group_464 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(464), clk => clk, reset => reset); --
    end block;
    -- CP-element group 465:  transition  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (6) 
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_sample_completed_
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_update_start_
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/$exit
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Sample/ack
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/req
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1470_inst_ack_0, ack => convTranspose_CP_34_elements(465)); -- 
    req_3426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(465), ack => WPIPE_ConvTranspose_output_pipe_1470_inst_req_1); -- 
    -- CP-element group 466:  transition  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/$exit
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/WPIPE_ConvTranspose_output_pipe_1470_Update/ack
      -- 
    ack_3427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1470_inst_ack_1, ack => convTranspose_CP_34_elements(466)); -- 
    -- CP-element group 467:  branch  join  transition  place  output  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	422 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	468 
    -- CP-element group 467: 	469 
    -- CP-element group 467:  members (10) 
      -- CP-element group 467: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483__exit__
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484__entry__
      -- CP-element group 467: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_dead_link/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_eval_test/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_eval_test/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_eval_test/branch_req
      -- CP-element group 467: 	 branch_block_stmt_38/R_exitcond1_1485_place
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_if_link/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1484_else_link/$entry
      -- 
    branch_req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(467), ack => if_stmt_1484_branch_req_0); -- 
    convTranspose_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(422) & convTranspose_CP_34_elements(466);
      gj_convTranspose_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  merge  transition  place  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	467 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	497 
    -- CP-element group 468:  members (13) 
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490__exit__
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500
      -- CP-element group 468: 	 branch_block_stmt_38/if_stmt_1484_if_link/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/if_stmt_1484_if_link/if_choice_transition
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiReqMerge
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiAck/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiAck/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/merge_stmt_1490_PhiAck/dummy
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500_PhiReq/$exit
      -- 
    if_choice_transition_3440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1484_branch_ack_1, ack => convTranspose_CP_34_elements(468)); -- 
    -- CP-element group 469:  fork  transition  place  input  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	467 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	492 
    -- CP-element group 469: 	493 
    -- CP-element group 469:  members (12) 
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_1484_else_link/$exit
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_1484_else_link/else_choice_transition
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1484_branch_ack_0, ack => convTranspose_CP_34_elements(469)); -- 
    rr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(469), ack => type_cast_1362_inst_req_0); -- 
    cr_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(469), ack => type_cast_1362_inst_req_1); -- 
    -- CP-element group 470:  merge  branch  transition  place  output  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	120 
    -- CP-element group 470: 	165 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	121 
    -- CP-element group 470: 	122 
    -- CP-element group 470:  members (17) 
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429__exit__
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435__entry__
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435__exit__
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436__entry__
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/assign_stmt_435/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_dead_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_eval_test/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_eval_test/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_eval_test/branch_req
      -- CP-element group 470: 	 branch_block_stmt_38/R_cmp194509_437_place
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_if_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/if_stmt_436_else_link/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiReqMerge
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/$entry
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/dummy
      -- 
    branch_req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(470), ack => if_stmt_436_branch_req_0); -- 
    convTranspose_CP_34_elements(470) <= OrReduce(convTranspose_CP_34_elements(120) & convTranspose_CP_34_elements(165));
    -- CP-element group 471:  transition  output  delay-element  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	124 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	475 
    -- CP-element group 471:  members (5) 
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_478_konst_delay_trans
      -- CP-element group 471: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_req
      -- 
    phi_stmt_474_req_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_474_req_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(471), ack => phi_stmt_474_req_0); -- 
    -- Element group convTranspose_CP_34_elements(471) is a control-delay.
    cp_element_471_delay: control_delay_element  generic map(name => " 471_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(124), ack => convTranspose_CP_34_elements(471), clk => clk, reset =>reset);
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	166 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	474 
    -- CP-element group 472:  members (2) 
      -- CP-element group 472: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/ra
      -- 
    ra_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_0, ack => convTranspose_CP_34_elements(472)); -- 
    -- CP-element group 473:  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	166 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (2) 
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/ca
      -- 
    ca_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_1, ack => convTranspose_CP_34_elements(473)); -- 
    -- CP-element group 474:  join  transition  output  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	472 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (6) 
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/$exit
      -- CP-element group 474: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_req
      -- 
    phi_stmt_474_req_3518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_474_req_3518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(474), ack => phi_stmt_474_req_1); -- 
    convTranspose_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(472) & convTranspose_CP_34_elements(473);
      gj_convTranspose_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  merge  transition  place  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	471 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (2) 
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473_PhiReqMerge
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(475) <= OrReduce(convTranspose_CP_34_elements(471) & convTranspose_CP_34_elements(474));
    -- CP-element group 476:  fork  transition  place  input  output  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	125 
    -- CP-element group 476: 	126 
    -- CP-element group 476: 	128 
    -- CP-element group 476: 	129 
    -- CP-element group 476: 	132 
    -- CP-element group 476: 	136 
    -- CP-element group 476: 	140 
    -- CP-element group 476: 	144 
    -- CP-element group 476: 	148 
    -- CP-element group 476: 	152 
    -- CP-element group 476: 	156 
    -- CP-element group 476: 	160 
    -- CP-element group 476: 	163 
    -- CP-element group 476:  members (56) 
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/merge_stmt_473__exit__
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636__entry__
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resized_1
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scaled_1
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_computed_1
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/index_resize_req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/index_resize_ack
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/scale_rename_req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/scale_rename_ack
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_update_start
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/req
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_sample_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/rr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_update_start_
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/$entry
      -- CP-element group 476: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/cr
      -- CP-element group 476: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/phi_stmt_474_ack
      -- 
    phi_stmt_474_ack_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_474_ack_0, ack => convTranspose_CP_34_elements(476)); -- 
    cr_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_615_inst_req_1); -- 
    cr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_543_inst_req_1); -- 
    cr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => ptr_deref_623_store_0_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_579_inst_req_1); -- 
    cr_1140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_561_inst_req_1); -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_597_inst_req_1); -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => array_obj_ref_486_index_offset_req_0); -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => array_obj_ref_486_index_offset_req_1); -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => addr_of_487_final_reg_req_1); -- 
    rr_1009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => RPIPE_ConvTranspose_input_pipe_490_inst_req_0); -- 
    cr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_494_inst_req_1); -- 
    cr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_507_inst_req_1); -- 
    cr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => type_cast_525_inst_req_1); -- 
    -- CP-element group 477:  transition  output  delay-element  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	168 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	481 
    -- CP-element group 477:  members (5) 
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_685_konst_delay_trans
      -- CP-element group 477: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_req
      -- 
    phi_stmt_681_req_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_req_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(477), ack => phi_stmt_681_req_0); -- 
    -- Element group convTranspose_CP_34_elements(477) is a control-delay.
    cp_element_477_delay: control_delay_element  generic map(name => " 477_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(168), ack => convTranspose_CP_34_elements(477), clk => clk, reset =>reset);
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	210 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	480 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/$exit
      -- CP-element group 478: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/ra
      -- 
    ra_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_0, ack => convTranspose_CP_34_elements(478)); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	210 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (2) 
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/ca
      -- 
    ca_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_1, ack => convTranspose_CP_34_elements(479)); -- 
    -- CP-element group 480:  join  transition  output  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	478 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (6) 
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/$exit
      -- CP-element group 480: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_req
      -- 
    phi_stmt_681_req_3572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_req_3572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(480), ack => phi_stmt_681_req_1); -- 
    convTranspose_cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_480"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(478) & convTranspose_CP_34_elements(479);
      gj_convTranspose_cp_element_group_480 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481:  merge  transition  place  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	477 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481:  members (2) 
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680_PhiReqMerge
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(481) <= OrReduce(convTranspose_CP_34_elements(477) & convTranspose_CP_34_elements(480));
    -- CP-element group 482:  fork  transition  place  input  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	169 
    -- CP-element group 482: 	170 
    -- CP-element group 482: 	172 
    -- CP-element group 482: 	173 
    -- CP-element group 482: 	176 
    -- CP-element group 482: 	180 
    -- CP-element group 482: 	184 
    -- CP-element group 482: 	188 
    -- CP-element group 482: 	192 
    -- CP-element group 482: 	196 
    -- CP-element group 482: 	200 
    -- CP-element group 482: 	204 
    -- CP-element group 482: 	207 
    -- CP-element group 482:  members (56) 
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_680__exit__
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843__entry__
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_update_start
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/scale_rename_ack
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/scale_rename_req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/index_resize_ack
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/index_resize_req
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_computed_1
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scaled_1
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resized_1
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/cr
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/phi_stmt_681_ack
      -- 
    phi_stmt_681_ack_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_681_ack_0, ack => convTranspose_CP_34_elements(482)); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => array_obj_ref_693_index_offset_req_1); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => array_obj_ref_693_index_offset_req_0); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_714_inst_req_1); -- 
    cr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_732_inst_req_1); -- 
    rr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => RPIPE_ConvTranspose_input_pipe_697_inst_req_0); -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => addr_of_694_final_reg_req_1); -- 
    cr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_701_inst_req_1); -- 
    cr_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_750_inst_req_1); -- 
    cr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_768_inst_req_1); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_786_inst_req_1); -- 
    cr_1555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_804_inst_req_1); -- 
    cr_1583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_822_inst_req_1); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => ptr_deref_830_store_0_req_1); -- 
    -- CP-element group 483:  merge  fork  transition  place  output  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	122 
    -- CP-element group 483: 	209 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	213 
    -- CP-element group 483: 	214 
    -- CP-element group 483: 	215 
    -- CP-element group 483: 	216 
    -- CP-element group 483: 	211 
    -- CP-element group 483: 	212 
    -- CP-element group 483:  members (25) 
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852__exit__
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880__entry__
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_update_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/cr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_update_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/cr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_sample_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_update_start_
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/rr
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/cr
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiReqMerge
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/$entry
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/$exit
      -- CP-element group 483: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/dummy
      -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_855_inst_req_0); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_855_inst_req_1); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_859_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_859_inst_req_1); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_863_inst_req_0); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => type_cast_863_inst_req_1); -- 
    convTranspose_CP_34_elements(483) <= OrReduce(convTranspose_CP_34_elements(122) & convTranspose_CP_34_elements(209));
    -- CP-element group 484:  transition  output  delay-element  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	221 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	488 
    -- CP-element group 484:  members (5) 
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_931_konst_delay_trans
      -- CP-element group 484: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_req
      -- 
    phi_stmt_925_req_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_925_req_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(484), ack => phi_stmt_925_req_1); -- 
    -- Element group convTranspose_CP_34_elements(484) is a control-delay.
    cp_element_484_delay: control_delay_element  generic map(name => " 484_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(221), ack => convTranspose_CP_34_elements(484), clk => clk, reset =>reset);
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	230 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	487 
    -- CP-element group 485:  members (2) 
      -- CP-element group 485: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/ra
      -- 
    ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_0, ack => convTranspose_CP_34_elements(485)); -- 
    -- CP-element group 486:  transition  input  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	230 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (2) 
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/ca
      -- 
    ca_3648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_1, ack => convTranspose_CP_34_elements(486)); -- 
    -- CP-element group 487:  join  transition  output  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	485 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (6) 
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/$exit
      -- CP-element group 487: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_req
      -- 
    phi_stmt_925_req_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_925_req_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(487), ack => phi_stmt_925_req_0); -- 
    convTranspose_cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_487"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(485) & convTranspose_CP_34_elements(486);
      gj_convTranspose_cp_element_group_487 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(487), clk => clk, reset => reset); --
    end block;
    -- CP-element group 488:  merge  transition  place  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	484 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (2) 
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924_PhiReqMerge
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(488) <= OrReduce(convTranspose_CP_34_elements(484) & convTranspose_CP_34_elements(487));
    -- CP-element group 489:  fork  transition  place  input  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	222 
    -- CP-element group 489: 	223 
    -- CP-element group 489: 	225 
    -- CP-element group 489: 	227 
    -- CP-element group 489:  members (29) 
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_924__exit__
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955__entry__
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_update_start_
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resized_1
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scaled_1
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_computed_1
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/index_resize_req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/index_resize_ack
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/scale_rename_req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/scale_rename_ack
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_update_start
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/req
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_update_start_
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/cr
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/phi_stmt_925_ack
      -- 
    phi_stmt_925_ack_3654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_925_ack_0, ack => convTranspose_CP_34_elements(489)); -- 
    req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => array_obj_ref_937_index_offset_req_0); -- 
    req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => array_obj_ref_937_index_offset_req_1); -- 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => addr_of_938_final_reg_req_1); -- 
    cr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => ptr_deref_941_store_0_req_1); -- 
    -- CP-element group 490:  merge  fork  transition  place  output  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	219 
    -- CP-element group 490: 	229 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	231 
    -- CP-element group 490: 	232 
    -- CP-element group 490: 	234 
    -- CP-element group 490:  members (16) 
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964__exit__
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973__entry__
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_update_start_
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/crr
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/ccr
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_update_start_
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/cr
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiReqMerge
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/$entry
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/$exit
      -- CP-element group 490: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/dummy
      -- 
    crr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => call_stmt_967_call_req_0); -- 
    ccr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => call_stmt_967_call_req_1); -- 
    cr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => type_cast_972_inst_req_1); -- 
    convTranspose_CP_34_elements(490) <= OrReduce(convTranspose_CP_34_elements(219) & convTranspose_CP_34_elements(229));
    -- CP-element group 491:  transition  output  delay-element  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	421 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	495 
    -- CP-element group 491:  members (5) 
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1360_konst_delay_trans
      -- CP-element group 491: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_req
      -- 
    phi_stmt_1356_req_3700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1356_req_3700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(491), ack => phi_stmt_1356_req_0); -- 
    -- Element group convTranspose_CP_34_elements(491) is a control-delay.
    cp_element_491_delay: control_delay_element  generic map(name => " 491_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(421), ack => convTranspose_CP_34_elements(491), clk => clk, reset =>reset);
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	469 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	494 
    -- CP-element group 492:  members (2) 
      -- CP-element group 492: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/$exit
      -- CP-element group 492: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Sample/ra
      -- 
    ra_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1362_inst_ack_0, ack => convTranspose_CP_34_elements(492)); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	469 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (2) 
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/Update/ca
      -- 
    ca_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1362_inst_ack_1, ack => convTranspose_CP_34_elements(493)); -- 
    -- CP-element group 494:  join  transition  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	492 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (6) 
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_sources/type_cast_1362/SplitProtocol/$exit
      -- CP-element group 494: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1356/phi_stmt_1356_req
      -- 
    phi_stmt_1356_req_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1356_req_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(494), ack => phi_stmt_1356_req_1); -- 
    convTranspose_cp_element_group_494: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_494"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(492) & convTranspose_CP_34_elements(493);
      gj_convTranspose_cp_element_group_494 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(494), clk => clk, reset => reset); --
    end block;
    -- CP-element group 495:  merge  transition  place  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	491 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (2) 
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1355_PhiReqMerge
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1355_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(495) <= OrReduce(convTranspose_CP_34_elements(491) & convTranspose_CP_34_elements(494));
    -- CP-element group 496:  fork  transition  place  input  output  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	422 
    -- CP-element group 496: 	423 
    -- CP-element group 496: 	425 
    -- CP-element group 496: 	427 
    -- CP-element group 496: 	429 
    -- CP-element group 496: 	431 
    -- CP-element group 496: 	433 
    -- CP-element group 496: 	435 
    -- CP-element group 496: 	437 
    -- CP-element group 496: 	439 
    -- CP-element group 496: 	441 
    -- CP-element group 496: 	443 
    -- CP-element group 496:  members (53) 
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1355__exit__
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483__entry__
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/word_0/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/scale_rename_req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1417_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/index_resize_req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/word_access_complete/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resized_1
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scaled_1
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_resize_1/index_resize_ack
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_computed_1
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_index_scale_1/scale_rename_ack
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1387_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1377_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1407_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/ptr_deref_1373_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/addr_of_1369_complete/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1427_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1447_update_start_
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/cr
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1397_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/req
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/type_cast_1437_Update/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_Sample/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/assign_stmt_1370_to_assign_stmt_1483/array_obj_ref_1368_final_index_sum_regn_update_start
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1355_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1355_PhiAck/phi_stmt_1356_ack
      -- 
    phi_stmt_1356_ack_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1356_ack_0, ack => convTranspose_CP_34_elements(496)); -- 
    cr_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => ptr_deref_1373_load_0_req_1); -- 
    cr_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1417_inst_req_1); -- 
    cr_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1387_inst_req_1); -- 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1427_inst_req_1); -- 
    cr_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1377_inst_req_1); -- 
    cr_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1407_inst_req_1); -- 
    req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => addr_of_1369_final_reg_req_1); -- 
    cr_3314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1447_inst_req_1); -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1397_inst_req_1); -- 
    req_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => array_obj_ref_1368_index_offset_req_1); -- 
    cr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => type_cast_1437_inst_req_1); -- 
    req_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(496), ack => array_obj_ref_1368_index_offset_req_0); -- 
    -- CP-element group 497:  merge  transition  place  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	419 
    -- CP-element group 497: 	468 
    -- CP-element group 497: successors 
    -- CP-element group 497:  members (16) 
      -- CP-element group 497: 	 $exit
      -- CP-element group 497: 	 branch_block_stmt_38/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/branch_block_stmt_38__exit__
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492__exit__
      -- CP-element group 497: 	 branch_block_stmt_38/return__
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494__exit__
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiReqMerge
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiAck/$entry
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiAck/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1492_PhiAck/dummy
      -- CP-element group 497: 	 branch_block_stmt_38/return___PhiReq/$entry
      -- CP-element group 497: 	 branch_block_stmt_38/return___PhiReq/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiReqMerge
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiAck/$entry
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiAck/$exit
      -- CP-element group 497: 	 branch_block_stmt_38/merge_stmt_1494_PhiAck/dummy
      -- 
    convTranspose_CP_34_elements(497) <= OrReduce(convTranspose_CP_34_elements(419) & convTranspose_CP_34_elements(468));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar525_936_resized : std_logic_vector(13 downto 0);
    signal R_indvar525_936_scaled : std_logic_vector(13 downto 0);
    signal R_indvar539_692_resized : std_logic_vector(10 downto 0);
    signal R_indvar539_692_scaled : std_logic_vector(10 downto 0);
    signal R_indvar555_485_resized : std_logic_vector(13 downto 0);
    signal R_indvar555_485_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1367_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1367_scaled : std_logic_vector(13 downto 0);
    signal add108_339 : std_logic_vector(15 downto 0);
    signal add117_364 : std_logic_vector(15 downto 0);
    signal add126_389 : std_logic_vector(15 downto 0);
    signal add12_88 : std_logic_vector(15 downto 0);
    signal add135_414 : std_logic_vector(15 downto 0);
    signal add150_513 : std_logic_vector(63 downto 0);
    signal add156_531 : std_logic_vector(63 downto 0);
    signal add162_549 : std_logic_vector(63 downto 0);
    signal add168_567 : std_logic_vector(63 downto 0);
    signal add174_585 : std_logic_vector(63 downto 0);
    signal add180_603 : std_logic_vector(63 downto 0);
    signal add186_621 : std_logic_vector(63 downto 0);
    signal add206_720 : std_logic_vector(63 downto 0);
    signal add212_738 : std_logic_vector(63 downto 0);
    signal add218_756 : std_logic_vector(63 downto 0);
    signal add21_113 : std_logic_vector(15 downto 0);
    signal add224_774 : std_logic_vector(63 downto 0);
    signal add230_792 : std_logic_vector(63 downto 0);
    signal add236_810 : std_logic_vector(63 downto 0);
    signal add242_828 : std_logic_vector(63 downto 0);
    signal add30_138 : std_logic_vector(15 downto 0);
    signal add39_163 : std_logic_vector(15 downto 0);
    signal add48_188 : std_logic_vector(15 downto 0);
    signal add57_213 : std_logic_vector(15 downto 0);
    signal add74_253 : std_logic_vector(31 downto 0);
    signal add79_258 : std_logic_vector(31 downto 0);
    signal add99_314 : std_logic_vector(15 downto 0);
    signal add_63 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1368_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1368_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_693_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_937_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_695 : std_logic_vector(31 downto 0);
    signal arrayidx269_939 : std_logic_vector(31 downto 0);
    signal arrayidx432_1370 : std_logic_vector(31 downto 0);
    signal arrayidx_488 : std_logic_vector(31 downto 0);
    signal call101_317 : std_logic_vector(7 downto 0);
    signal call106_330 : std_logic_vector(7 downto 0);
    signal call10_79 : std_logic_vector(7 downto 0);
    signal call110_342 : std_logic_vector(7 downto 0);
    signal call115_355 : std_logic_vector(7 downto 0);
    signal call119_367 : std_logic_vector(7 downto 0);
    signal call124_380 : std_logic_vector(7 downto 0);
    signal call128_392 : std_logic_vector(7 downto 0);
    signal call133_405 : std_logic_vector(7 downto 0);
    signal call143_491 : std_logic_vector(7 downto 0);
    signal call147_504 : std_logic_vector(7 downto 0);
    signal call14_91 : std_logic_vector(7 downto 0);
    signal call153_522 : std_logic_vector(7 downto 0);
    signal call159_540 : std_logic_vector(7 downto 0);
    signal call165_558 : std_logic_vector(7 downto 0);
    signal call171_576 : std_logic_vector(7 downto 0);
    signal call177_594 : std_logic_vector(7 downto 0);
    signal call183_612 : std_logic_vector(7 downto 0);
    signal call199_698 : std_logic_vector(7 downto 0);
    signal call19_104 : std_logic_vector(7 downto 0);
    signal call203_711 : std_logic_vector(7 downto 0);
    signal call209_729 : std_logic_vector(7 downto 0);
    signal call215_747 : std_logic_vector(7 downto 0);
    signal call221_765 : std_logic_vector(7 downto 0);
    signal call227_783 : std_logic_vector(7 downto 0);
    signal call233_801 : std_logic_vector(7 downto 0);
    signal call239_819 : std_logic_vector(7 downto 0);
    signal call23_116 : std_logic_vector(7 downto 0);
    signal call275_967 : std_logic_vector(63 downto 0);
    signal call28_129 : std_logic_vector(7 downto 0);
    signal call2_54 : std_logic_vector(7 downto 0);
    signal call32_141 : std_logic_vector(7 downto 0);
    signal call346_1190 : std_logic_vector(15 downto 0);
    signal call348_1193 : std_logic_vector(15 downto 0);
    signal call350_1196 : std_logic_vector(15 downto 0);
    signal call352_1199 : std_logic_vector(15 downto 0);
    signal call354_1202 : std_logic_vector(63 downto 0);
    signal call37_154 : std_logic_vector(7 downto 0);
    signal call41_166 : std_logic_vector(7 downto 0);
    signal call46_179 : std_logic_vector(7 downto 0);
    signal call50_191 : std_logic_vector(7 downto 0);
    signal call55_204 : std_logic_vector(7 downto 0);
    signal call5_66 : std_logic_vector(7 downto 0);
    signal call92_292 : std_logic_vector(7 downto 0);
    signal call97_305 : std_logic_vector(7 downto 0);
    signal call_41 : std_logic_vector(7 downto 0);
    signal cmp194509_435 : std_logic_vector(0 downto 0);
    signal cmp264505_880 : std_logic_vector(0 downto 0);
    signal cmp513_420 : std_logic_vector(0 downto 0);
    signal conv104_321 : std_logic_vector(15 downto 0);
    signal conv107_334 : std_logic_vector(15 downto 0);
    signal conv113_346 : std_logic_vector(15 downto 0);
    signal conv116_359 : std_logic_vector(15 downto 0);
    signal conv11_83 : std_logic_vector(15 downto 0);
    signal conv122_371 : std_logic_vector(15 downto 0);
    signal conv125_384 : std_logic_vector(15 downto 0);
    signal conv131_396 : std_logic_vector(15 downto 0);
    signal conv134_409 : std_logic_vector(15 downto 0);
    signal conv144_495 : std_logic_vector(63 downto 0);
    signal conv149_508 : std_logic_vector(63 downto 0);
    signal conv155_526 : std_logic_vector(63 downto 0);
    signal conv161_544 : std_logic_vector(63 downto 0);
    signal conv167_562 : std_logic_vector(63 downto 0);
    signal conv173_580 : std_logic_vector(63 downto 0);
    signal conv179_598 : std_logic_vector(63 downto 0);
    signal conv17_95 : std_logic_vector(15 downto 0);
    signal conv185_616 : std_logic_vector(63 downto 0);
    signal conv1_45 : std_logic_vector(15 downto 0);
    signal conv200_702 : std_logic_vector(63 downto 0);
    signal conv205_715 : std_logic_vector(63 downto 0);
    signal conv20_108 : std_logic_vector(15 downto 0);
    signal conv211_733 : std_logic_vector(63 downto 0);
    signal conv217_751 : std_logic_vector(63 downto 0);
    signal conv223_769 : std_logic_vector(63 downto 0);
    signal conv229_787 : std_logic_vector(63 downto 0);
    signal conv235_805 : std_logic_vector(63 downto 0);
    signal conv241_823 : std_logic_vector(63 downto 0);
    signal conv253_856 : std_logic_vector(31 downto 0);
    signal conv255_860 : std_logic_vector(31 downto 0);
    signal conv258_864 : std_logic_vector(31 downto 0);
    signal conv26_120 : std_logic_vector(15 downto 0);
    signal conv276_973 : std_logic_vector(63 downto 0);
    signal conv29_133 : std_logic_vector(15 downto 0);
    signal conv305_1055 : std_logic_vector(15 downto 0);
    signal conv307_1062 : std_logic_vector(15 downto 0);
    signal conv322_1111 : std_logic_vector(15 downto 0);
    signal conv324_1118 : std_logic_vector(15 downto 0);
    signal conv339_1167 : std_logic_vector(15 downto 0);
    signal conv341_1174 : std_logic_vector(15 downto 0);
    signal conv355_1207 : std_logic_vector(63 downto 0);
    signal conv35_145 : std_logic_vector(15 downto 0);
    signal conv361_1216 : std_logic_vector(7 downto 0);
    signal conv367_1226 : std_logic_vector(7 downto 0);
    signal conv373_1236 : std_logic_vector(7 downto 0);
    signal conv379_1246 : std_logic_vector(7 downto 0);
    signal conv385_1256 : std_logic_vector(7 downto 0);
    signal conv38_158 : std_logic_vector(15 downto 0);
    signal conv391_1266 : std_logic_vector(7 downto 0);
    signal conv397_1276 : std_logic_vector(7 downto 0);
    signal conv3_58 : std_logic_vector(15 downto 0);
    signal conv403_1286 : std_logic_vector(7 downto 0);
    signal conv437_1378 : std_logic_vector(7 downto 0);
    signal conv443_1388 : std_logic_vector(7 downto 0);
    signal conv449_1398 : std_logic_vector(7 downto 0);
    signal conv44_170 : std_logic_vector(15 downto 0);
    signal conv455_1408 : std_logic_vector(7 downto 0);
    signal conv461_1418 : std_logic_vector(7 downto 0);
    signal conv467_1428 : std_logic_vector(7 downto 0);
    signal conv473_1438 : std_logic_vector(7 downto 0);
    signal conv479_1448 : std_logic_vector(7 downto 0);
    signal conv47_183 : std_logic_vector(15 downto 0);
    signal conv53_195 : std_logic_vector(15 downto 0);
    signal conv56_208 : std_logic_vector(15 downto 0);
    signal conv61_217 : std_logic_vector(31 downto 0);
    signal conv63_221 : std_logic_vector(31 downto 0);
    signal conv65_225 : std_logic_vector(31 downto 0);
    signal conv82_262 : std_logic_vector(31 downto 0);
    signal conv84_266 : std_logic_vector(31 downto 0);
    signal conv87_270 : std_logic_vector(31 downto 0);
    signal conv8_70 : std_logic_vector(15 downto 0);
    signal conv90_274 : std_logic_vector(31 downto 0);
    signal conv95_296 : std_logic_vector(15 downto 0);
    signal conv98_309 : std_logic_vector(15 downto 0);
    signal exitcond1_1483 : std_logic_vector(0 downto 0);
    signal exitcond2_843 : std_logic_vector(0 downto 0);
    signal exitcond3_636 : std_logic_vector(0 downto 0);
    signal exitcond_955 : std_logic_vector(0 downto 0);
    signal iNsTr_14_247 : std_logic_vector(31 downto 0);
    signal iNsTr_196_1340 : std_logic_vector(63 downto 0);
    signal iNsTr_26_458 : std_logic_vector(63 downto 0);
    signal iNsTr_39_665 : std_logic_vector(63 downto 0);
    signal iNsTr_53_909 : std_logic_vector(63 downto 0);
    signal indvar525_925 : std_logic_vector(63 downto 0);
    signal indvar539_681 : std_logic_vector(63 downto 0);
    signal indvar555_474 : std_logic_vector(63 downto 0);
    signal indvar_1356 : std_logic_vector(63 downto 0);
    signal indvarx_xnext526_950 : std_logic_vector(63 downto 0);
    signal indvarx_xnext540_838 : std_logic_vector(63 downto 0);
    signal indvarx_xnext556_631 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1478 : std_logic_vector(63 downto 0);
    signal mul256_869 : std_logic_vector(31 downto 0);
    signal mul259_874 : std_logic_vector(31 downto 0);
    signal mul66_235 : std_logic_vector(31 downto 0);
    signal mul85_279 : std_logic_vector(31 downto 0);
    signal mul88_284 : std_logic_vector(31 downto 0);
    signal mul91_289 : std_logic_vector(31 downto 0);
    signal mul_230 : std_logic_vector(31 downto 0);
    signal ptr_deref_1373_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1373_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1373_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1373_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1373_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_623_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_623_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_623_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_623_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_623_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_623_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_830_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_830_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_830_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_830_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_830_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_830_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_941_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_941_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_941_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_941_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_941_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_941_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_327 : std_logic_vector(15 downto 0);
    signal shl114_352 : std_logic_vector(15 downto 0);
    signal shl123_377 : std_logic_vector(15 downto 0);
    signal shl132_402 : std_logic_vector(15 downto 0);
    signal shl146_501 : std_logic_vector(63 downto 0);
    signal shl152_519 : std_logic_vector(63 downto 0);
    signal shl158_537 : std_logic_vector(63 downto 0);
    signal shl164_555 : std_logic_vector(63 downto 0);
    signal shl170_573 : std_logic_vector(63 downto 0);
    signal shl176_591 : std_logic_vector(63 downto 0);
    signal shl182_609 : std_logic_vector(63 downto 0);
    signal shl18_101 : std_logic_vector(15 downto 0);
    signal shl202_708 : std_logic_vector(63 downto 0);
    signal shl208_726 : std_logic_vector(63 downto 0);
    signal shl214_744 : std_logic_vector(63 downto 0);
    signal shl220_762 : std_logic_vector(63 downto 0);
    signal shl226_780 : std_logic_vector(63 downto 0);
    signal shl232_798 : std_logic_vector(63 downto 0);
    signal shl238_816 : std_logic_vector(63 downto 0);
    signal shl27_126 : std_logic_vector(15 downto 0);
    signal shl36_151 : std_logic_vector(15 downto 0);
    signal shl45_176 : std_logic_vector(15 downto 0);
    signal shl54_201 : std_logic_vector(15 downto 0);
    signal shl96_302 : std_logic_vector(15 downto 0);
    signal shl9_76 : std_logic_vector(15 downto 0);
    signal shl_51 : std_logic_vector(15 downto 0);
    signal shr304_1051 : std_logic_vector(31 downto 0);
    signal shr321_1107 : std_logic_vector(31 downto 0);
    signal shr338_1163 : std_logic_vector(31 downto 0);
    signal shr364_1222 : std_logic_vector(63 downto 0);
    signal shr370_1232 : std_logic_vector(63 downto 0);
    signal shr376_1242 : std_logic_vector(63 downto 0);
    signal shr382_1252 : std_logic_vector(63 downto 0);
    signal shr388_1262 : std_logic_vector(63 downto 0);
    signal shr394_1272 : std_logic_vector(63 downto 0);
    signal shr400_1282 : std_logic_vector(63 downto 0);
    signal shr440_1384 : std_logic_vector(63 downto 0);
    signal shr446_1394 : std_logic_vector(63 downto 0);
    signal shr452_1404 : std_logic_vector(63 downto 0);
    signal shr458_1414 : std_logic_vector(63 downto 0);
    signal shr464_1424 : std_logic_vector(63 downto 0);
    signal shr470_1434 : std_logic_vector(63 downto 0);
    signal shr476_1444 : std_logic_vector(63 downto 0);
    signal shr_241 : std_logic_vector(31 downto 0);
    signal sub_1212 : std_logic_vector(63 downto 0);
    signal tmp433_1374 : std_logic_vector(63 downto 0);
    signal tmp520_1324 : std_logic_vector(31 downto 0);
    signal tmp520x_xop_1336 : std_logic_vector(31 downto 0);
    signal tmp521_1330 : std_logic_vector(0 downto 0);
    signal tmp524_1353 : std_logic_vector(63 downto 0);
    signal tmp532_893 : std_logic_vector(31 downto 0);
    signal tmp532x_xop_905 : std_logic_vector(31 downto 0);
    signal tmp533_899 : std_logic_vector(0 downto 0);
    signal tmp537_922 : std_logic_vector(63 downto 0);
    signal tmp548_649 : std_logic_vector(31 downto 0);
    signal tmp548x_xop_661 : std_logic_vector(31 downto 0);
    signal tmp549_655 : std_logic_vector(0 downto 0);
    signal tmp553_678 : std_logic_vector(63 downto 0);
    signal tmp562x_xop_454 : std_logic_vector(31 downto 0);
    signal tmp563_448 : std_logic_vector(0 downto 0);
    signal tmp567_471 : std_logic_vector(63 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1161_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1205_wire : std_logic_vector(63 downto 0);
    signal type_cast_1220_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1230_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1240_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_124_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1250_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1270_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1280_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1328_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1360_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1362_wire : std_logic_vector(63 downto 0);
    signal type_cast_1382_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1392_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1402_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1412_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1442_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1476_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_149_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_174_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_300_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_375_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_400_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_418_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_462_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_469_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_480_wire : std_logic_vector(63 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_517_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_535_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_571_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_589_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_629_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_653_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_659_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_669_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_685_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_687_wire : std_logic_vector(63 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_742_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_74_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_814_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_928_wire : std_logic_vector(63 downto 0);
    signal type_cast_931_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_971_wire : std_logic_vector(63 downto 0);
    signal type_cast_99_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop569_915 : std_logic_vector(63 downto 0);
    signal xx_xop570_671 : std_logic_vector(63 downto 0);
    signal xx_xop571_464 : std_logic_vector(63 downto 0);
    signal xx_xop_1346 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1368_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1368_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1368_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1368_resized_base_address <= "00000000000000";
    array_obj_ref_486_constant_part_of_offset <= "00000000000000";
    array_obj_ref_486_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_486_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_486_resized_base_address <= "00000000000000";
    array_obj_ref_693_constant_part_of_offset <= "00000100010";
    array_obj_ref_693_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_693_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_693_resized_base_address <= "00000000000";
    array_obj_ref_937_constant_part_of_offset <= "00000000000000";
    array_obj_ref_937_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_937_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_937_resized_base_address <= "00000000000000";
    ptr_deref_1373_word_offset_0 <= "00000000000000";
    ptr_deref_623_word_offset_0 <= "00000000000000";
    ptr_deref_830_word_offset_0 <= "00000000000";
    ptr_deref_941_word_offset_0 <= "00000000000000";
    type_cast_1004_wire_constant <= "0000000000000000";
    type_cast_1008_wire_constant <= "0000000000000000";
    type_cast_1049_wire_constant <= "00000000000000000000000000010010";
    type_cast_1105_wire_constant <= "00000000000000000000000000010001";
    type_cast_1161_wire_constant <= "00000000000000000000000000010000";
    type_cast_1220_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1230_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1240_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_124_wire_constant <= "0000000000001000";
    type_cast_1250_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1260_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1270_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1280_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1322_wire_constant <= "00000000000000000000000000000010";
    type_cast_1328_wire_constant <= "00000000000000000000000000000001";
    type_cast_1334_wire_constant <= "11111111111111111111111111111111";
    type_cast_1344_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1351_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1360_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1382_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1392_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1402_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1412_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1432_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1442_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1476_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_149_wire_constant <= "0000000000001000";
    type_cast_174_wire_constant <= "0000000000001000";
    type_cast_199_wire_constant <= "0000000000001000";
    type_cast_239_wire_constant <= "00000000000000000000000000000010";
    type_cast_245_wire_constant <= "00000000000000000000000000000001";
    type_cast_251_wire_constant <= "01111111111111111111111111111110";
    type_cast_300_wire_constant <= "0000000000001000";
    type_cast_325_wire_constant <= "0000000000001000";
    type_cast_350_wire_constant <= "0000000000001000";
    type_cast_375_wire_constant <= "0000000000001000";
    type_cast_400_wire_constant <= "0000000000001000";
    type_cast_418_wire_constant <= "00000000000000000000000000000011";
    type_cast_433_wire_constant <= "00000000000000000000000000000011";
    type_cast_446_wire_constant <= "00000000000000000000000000000001";
    type_cast_452_wire_constant <= "11111111111111111111111111111111";
    type_cast_462_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_49_wire_constant <= "0000000000001000";
    type_cast_517_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_553_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_589_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_629_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_647_wire_constant <= "00000000000000000000000000000010";
    type_cast_653_wire_constant <= "00000000000000000000000000000001";
    type_cast_659_wire_constant <= "11111111111111111111111111111111";
    type_cast_669_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_676_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_685_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_706_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_742_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_74_wire_constant <= "0000000000001000";
    type_cast_760_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_778_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_796_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_836_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_878_wire_constant <= "00000000000000000000000000000011";
    type_cast_891_wire_constant <= "00000000000000000000000000000010";
    type_cast_897_wire_constant <= "00000000000000000000000000000001";
    type_cast_903_wire_constant <= "11111111111111111111111111111111";
    type_cast_913_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_931_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_948_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_99_wire_constant <= "0000000000001000";
    phi_stmt_1356: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1360_wire_constant & type_cast_1362_wire;
      req <= phi_stmt_1356_req_0 & phi_stmt_1356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1356",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1356_ack_0,
          idata => idata,
          odata => indvar_1356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1356
    phi_stmt_474: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_478_wire_constant & type_cast_480_wire;
      req <= phi_stmt_474_req_0 & phi_stmt_474_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_474",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_474_ack_0,
          idata => idata,
          odata => indvar555_474,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_474
    phi_stmt_681: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_685_wire_constant & type_cast_687_wire;
      req <= phi_stmt_681_req_0 & phi_stmt_681_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_681",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_681_ack_0,
          idata => idata,
          odata => indvar539_681,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_681
    phi_stmt_925: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_928_wire & type_cast_931_wire_constant;
      req <= phi_stmt_925_req_0 & phi_stmt_925_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_925",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_925_ack_0,
          idata => idata,
          odata => indvar525_925,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_925
    -- flow-through select operator MUX_1352_inst
    tmp524_1353 <= xx_xop_1346 when (tmp521_1330(0) /=  '0') else type_cast_1351_wire_constant;
    -- flow-through select operator MUX_470_inst
    tmp567_471 <= xx_xop571_464 when (tmp563_448(0) /=  '0') else type_cast_469_wire_constant;
    -- flow-through select operator MUX_677_inst
    tmp553_678 <= xx_xop570_671 when (tmp549_655(0) /=  '0') else type_cast_676_wire_constant;
    -- flow-through select operator MUX_921_inst
    tmp537_922 <= xx_xop569_915 when (tmp533_899(0) /=  '0') else type_cast_920_wire_constant;
    addr_of_1369_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1369_final_reg_req_0;
      addr_of_1369_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1369_final_reg_req_1;
      addr_of_1369_final_reg_ack_1<= rack(0);
      addr_of_1369_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1369_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1368_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx432_1370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_487_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_487_final_reg_req_0;
      addr_of_487_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_487_final_reg_req_1;
      addr_of_487_final_reg_ack_1<= rack(0);
      addr_of_487_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_487_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_486_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_694_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_694_final_reg_req_0;
      addr_of_694_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_694_final_reg_req_1;
      addr_of_694_final_reg_ack_1<= rack(0);
      addr_of_694_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_694_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_693_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_938_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_938_final_reg_req_0;
      addr_of_938_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_938_final_reg_req_1;
      addr_of_938_final_reg_ack_1<= rack(0);
      addr_of_938_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_938_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_937_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_939,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1054_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1054_inst_req_0;
      type_cast_1054_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1054_inst_req_1;
      type_cast_1054_inst_ack_1<= rack(0);
      type_cast_1054_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1054_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1051,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1055,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1061_inst_req_0;
      type_cast_1061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1061_inst_req_1;
      type_cast_1061_inst_ack_1<= rack(0);
      type_cast_1061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_107_inst_req_0;
      type_cast_107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_107_inst_req_1;
      type_cast_107_inst_ack_1<= rack(0);
      type_cast_107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1117_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1117_inst_req_0;
      type_cast_1117_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1117_inst_req_1;
      type_cast_1117_inst_ack_1<= rack(0);
      type_cast_1117_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1117_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1166_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1166_inst_req_0;
      type_cast_1166_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1166_inst_req_1;
      type_cast_1166_inst_ack_1<= rack(0);
      type_cast_1166_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1166_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_119_inst_req_0;
      type_cast_119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_119_inst_req_1;
      type_cast_119_inst_ack_1<= rack(0);
      type_cast_119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1206_inst_req_0;
      type_cast_1206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1206_inst_req_1;
      type_cast_1206_inst_ack_1<= rack(0);
      type_cast_1206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1205_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1215_inst_req_0;
      type_cast_1215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1215_inst_req_1;
      type_cast_1215_inst_ack_1<= rack(0);
      type_cast_1215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv361_1216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1225_inst_req_0;
      type_cast_1225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1225_inst_req_1;
      type_cast_1225_inst_ack_1<= rack(0);
      type_cast_1225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr364_1222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1235_inst_req_0;
      type_cast_1235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1235_inst_req_1;
      type_cast_1235_inst_ack_1<= rack(0);
      type_cast_1235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr370_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1245_inst_req_0;
      type_cast_1245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1245_inst_req_1;
      type_cast_1245_inst_ack_1<= rack(0);
      type_cast_1245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr376_1242,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv379_1246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1255_inst_req_0;
      type_cast_1255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1255_inst_req_1;
      type_cast_1255_inst_ack_1<= rack(0);
      type_cast_1255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr382_1252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv385_1256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1265_inst_req_0;
      type_cast_1265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1265_inst_req_1;
      type_cast_1265_inst_ack_1<= rack(0);
      type_cast_1265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr388_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv391_1266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1275_inst_req_0;
      type_cast_1275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1275_inst_req_1;
      type_cast_1275_inst_ack_1<= rack(0);
      type_cast_1275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr394_1272,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv397_1276,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1285_inst_req_0;
      type_cast_1285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1285_inst_req_1;
      type_cast_1285_inst_ack_1<= rack(0);
      type_cast_1285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr400_1282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv403_1286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_132_inst_req_0;
      type_cast_132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_132_inst_req_1;
      type_cast_132_inst_ack_1<= rack(0);
      type_cast_132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1339_inst_req_0;
      type_cast_1339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1339_inst_req_1;
      type_cast_1339_inst_ack_1<= rack(0);
      type_cast_1339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp520x_xop_1336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_196_1340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1362_inst_req_0;
      type_cast_1362_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1362_inst_req_1;
      type_cast_1362_inst_ack_1<= rack(0);
      type_cast_1362_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1362_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1362_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1377_inst_req_0;
      type_cast_1377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1377_inst_req_1;
      type_cast_1377_inst_ack_1<= rack(0);
      type_cast_1377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp433_1374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv437_1378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1387_inst_req_0;
      type_cast_1387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1387_inst_req_1;
      type_cast_1387_inst_ack_1<= rack(0);
      type_cast_1387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr440_1384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv443_1388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1397_inst_req_0;
      type_cast_1397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1397_inst_req_1;
      type_cast_1397_inst_ack_1<= rack(0);
      type_cast_1397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr446_1394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv449_1398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1407_inst_req_0;
      type_cast_1407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1407_inst_req_1;
      type_cast_1407_inst_ack_1<= rack(0);
      type_cast_1407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr452_1404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv455_1408,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1417_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1417_inst_req_0;
      type_cast_1417_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1417_inst_req_1;
      type_cast_1417_inst_ack_1<= rack(0);
      type_cast_1417_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1417_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr458_1414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv461_1418,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1427_inst_req_0;
      type_cast_1427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1427_inst_req_1;
      type_cast_1427_inst_ack_1<= rack(0);
      type_cast_1427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr464_1424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv467_1428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1437_inst_req_0;
      type_cast_1437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1437_inst_req_1;
      type_cast_1437_inst_ack_1<= rack(0);
      type_cast_1437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr470_1434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv473_1438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1447_inst_req_0;
      type_cast_1447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1447_inst_req_1;
      type_cast_1447_inst_ack_1<= rack(0);
      type_cast_1447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr476_1444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1448,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_144_inst_req_0;
      type_cast_144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_144_inst_req_1;
      type_cast_144_inst_ack_1<= rack(0);
      type_cast_144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_157_inst_req_0;
      type_cast_157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_157_inst_req_1;
      type_cast_157_inst_ack_1<= rack(0);
      type_cast_157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_169_inst_req_0;
      type_cast_169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_169_inst_req_1;
      type_cast_169_inst_ack_1<= rack(0);
      type_cast_169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_166,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_207_inst_req_0;
      type_cast_207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_207_inst_req_1;
      type_cast_207_inst_ack_1<= rack(0);
      type_cast_207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_216_inst_req_0;
      type_cast_216_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_216_inst_req_1;
      type_cast_216_inst_ack_1<= rack(0);
      type_cast_216_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_216_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_220_inst_req_0;
      type_cast_220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_220_inst_req_1;
      type_cast_220_inst_ack_1<= rack(0);
      type_cast_220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_88,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_224_inst_req_0;
      type_cast_224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_224_inst_req_1;
      type_cast_224_inst_ack_1<= rack(0);
      type_cast_224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_261_inst_req_0;
      type_cast_261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_261_inst_req_1;
      type_cast_261_inst_ack_1<= rack(0);
      type_cast_261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_265_inst_req_0;
      type_cast_265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_265_inst_req_1;
      type_cast_265_inst_ack_1<= rack(0);
      type_cast_265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_273_inst_req_0;
      type_cast_273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_273_inst_req_1;
      type_cast_273_inst_ack_1<= rack(0);
      type_cast_273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_295_inst_req_0;
      type_cast_295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_295_inst_req_1;
      type_cast_295_inst_ack_1<= rack(0);
      type_cast_295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_308_inst_req_0;
      type_cast_308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_308_inst_req_1;
      type_cast_308_inst_ack_1<= rack(0);
      type_cast_308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_333_inst_req_0;
      type_cast_333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_333_inst_req_1;
      type_cast_333_inst_ack_1<= rack(0);
      type_cast_333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_383_inst_req_0;
      type_cast_383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_383_inst_req_1;
      type_cast_383_inst_ack_1<= rack(0);
      type_cast_383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_395_inst_req_0;
      type_cast_395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_395_inst_req_1;
      type_cast_395_inst_ack_1<= rack(0);
      type_cast_395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_408_inst_req_0;
      type_cast_408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_408_inst_req_1;
      type_cast_408_inst_ack_1<= rack(0);
      type_cast_408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_44_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_44_inst_req_0;
      type_cast_44_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_44_inst_req_1;
      type_cast_44_inst_ack_1<= rack(0);
      type_cast_44_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_44_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_45,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_457_inst_req_0;
      type_cast_457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_457_inst_req_1;
      type_cast_457_inst_ack_1<= rack(0);
      type_cast_457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp562x_xop_454,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_458,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_480_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_480_inst_req_0;
      type_cast_480_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_480_inst_req_1;
      type_cast_480_inst_ack_1<= rack(0);
      type_cast_480_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_480_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext556_631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_480_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_494_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_494_inst_req_0;
      type_cast_494_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_494_inst_req_1;
      type_cast_494_inst_ack_1<= rack(0);
      type_cast_494_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_494_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_491,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_507_inst_req_0;
      type_cast_507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_507_inst_req_1;
      type_cast_507_inst_ack_1<= rack(0);
      type_cast_507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_525_inst_req_0;
      type_cast_525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_525_inst_req_1;
      type_cast_525_inst_ack_1<= rack(0);
      type_cast_525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_543_inst_req_0;
      type_cast_543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_543_inst_req_1;
      type_cast_543_inst_ack_1<= rack(0);
      type_cast_543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_579_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_579_inst_req_0;
      type_cast_579_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_579_inst_req_1;
      type_cast_579_inst_ack_1<= rack(0);
      type_cast_579_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_579_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_576,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_580,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_57_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_57_inst_req_0;
      type_cast_57_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_57_inst_req_1;
      type_cast_57_inst_ack_1<= rack(0);
      type_cast_57_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_57_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_54,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_58,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_597_inst_req_0;
      type_cast_597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_597_inst_req_1;
      type_cast_597_inst_ack_1<= rack(0);
      type_cast_597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_615_inst_req_0;
      type_cast_615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_615_inst_req_1;
      type_cast_615_inst_ack_1<= rack(0);
      type_cast_615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_664_inst_req_0;
      type_cast_664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_664_inst_req_1;
      type_cast_664_inst_ack_1<= rack(0);
      type_cast_664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp548x_xop_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_687_inst_req_0;
      type_cast_687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_687_inst_req_1;
      type_cast_687_inst_ack_1<= rack(0);
      type_cast_687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext540_838,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_687_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_69_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_69_inst_req_0;
      type_cast_69_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_69_inst_req_1;
      type_cast_69_inst_ack_1<= rack(0);
      type_cast_69_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_69_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_66,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_70,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_701_inst_req_0;
      type_cast_701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_701_inst_req_1;
      type_cast_701_inst_ack_1<= rack(0);
      type_cast_701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_714_inst_req_0;
      type_cast_714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_714_inst_req_1;
      type_cast_714_inst_ack_1<= rack(0);
      type_cast_714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_732_inst_req_0;
      type_cast_732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_732_inst_req_1;
      type_cast_732_inst_ack_1<= rack(0);
      type_cast_732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_733,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_768_inst_req_0;
      type_cast_768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_768_inst_req_1;
      type_cast_768_inst_ack_1<= rack(0);
      type_cast_768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_786_inst_req_0;
      type_cast_786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_786_inst_req_1;
      type_cast_786_inst_ack_1<= rack(0);
      type_cast_786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_804_inst_req_0;
      type_cast_804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_804_inst_req_1;
      type_cast_804_inst_ack_1<= rack(0);
      type_cast_804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_805,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_822_inst_req_0;
      type_cast_822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_822_inst_req_1;
      type_cast_822_inst_ack_1<= rack(0);
      type_cast_822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_82_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_82_inst_req_0;
      type_cast_82_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_82_inst_req_1;
      type_cast_82_inst_ack_1<= rack(0);
      type_cast_82_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_82_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_79,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_83,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_855_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_855_inst_req_0;
      type_cast_855_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_855_inst_req_1;
      type_cast_855_inst_ack_1<= rack(0);
      type_cast_855_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_855_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_859_inst_req_0;
      type_cast_859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_859_inst_req_1;
      type_cast_859_inst_ack_1<= rack(0);
      type_cast_859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_863_inst_req_0;
      type_cast_863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_863_inst_req_1;
      type_cast_863_inst_ack_1<= rack(0);
      type_cast_863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_908_inst_req_0;
      type_cast_908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_908_inst_req_1;
      type_cast_908_inst_ack_1<= rack(0);
      type_cast_908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp532x_xop_905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_909,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_928_inst_req_0;
      type_cast_928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_928_inst_req_1;
      type_cast_928_inst_ack_1<= rack(0);
      type_cast_928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext526_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_928_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_94_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_94_inst_req_0;
      type_cast_94_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_94_inst_req_1;
      type_cast_94_inst_ack_1<= rack(0);
      type_cast_94_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_94_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_91,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_972_inst_req_0;
      type_cast_972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_972_inst_req_1;
      type_cast_972_inst_ack_1<= rack(0);
      type_cast_972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_971_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1368_index_1_rename
    process(R_indvar_1367_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1367_resized;
      ov(13 downto 0) := iv;
      R_indvar_1367_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1368_index_1_resize
    process(indvar_1356) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1356;
      ov := iv(13 downto 0);
      R_indvar_1367_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1368_root_address_inst
    process(array_obj_ref_1368_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1368_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1368_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_index_1_rename
    process(R_indvar555_485_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar555_485_resized;
      ov(13 downto 0) := iv;
      R_indvar555_485_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_index_1_resize
    process(indvar555_474) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar555_474;
      ov := iv(13 downto 0);
      R_indvar555_485_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_root_address_inst
    process(array_obj_ref_486_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_486_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_486_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_index_1_rename
    process(R_indvar539_692_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar539_692_resized;
      ov(10 downto 0) := iv;
      R_indvar539_692_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_index_1_resize
    process(indvar539_681) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar539_681;
      ov := iv(10 downto 0);
      R_indvar539_692_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_root_address_inst
    process(array_obj_ref_693_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_693_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_693_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_index_1_rename
    process(R_indvar525_936_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar525_936_resized;
      ov(13 downto 0) := iv;
      R_indvar525_936_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_index_1_resize
    process(indvar525_925) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar525_925;
      ov := iv(13 downto 0);
      R_indvar525_936_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_root_address_inst
    process(array_obj_ref_937_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_937_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_937_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_addr_0
    process(ptr_deref_1373_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1373_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1373_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_base_resize
    process(arrayidx432_1370) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx432_1370;
      ov := iv(13 downto 0);
      ptr_deref_1373_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_gather_scatter
    process(ptr_deref_1373_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1373_data_0;
      ov(63 downto 0) := iv;
      tmp433_1374 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1373_root_address_inst
    process(ptr_deref_1373_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1373_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1373_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_addr_0
    process(ptr_deref_623_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_623_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_623_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_base_resize
    process(arrayidx_488) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_488;
      ov := iv(13 downto 0);
      ptr_deref_623_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_gather_scatter
    process(add186_621) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_621;
      ov(63 downto 0) := iv;
      ptr_deref_623_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_root_address_inst
    process(ptr_deref_623_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_623_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_623_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_addr_0
    process(ptr_deref_830_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_830_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_830_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_base_resize
    process(arrayidx246_695) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_695;
      ov := iv(10 downto 0);
      ptr_deref_830_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_gather_scatter
    process(add242_828) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_828;
      ov(63 downto 0) := iv;
      ptr_deref_830_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_root_address_inst
    process(ptr_deref_830_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_830_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_830_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_addr_0
    process(ptr_deref_941_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_941_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_base_resize
    process(arrayidx269_939) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_939;
      ov := iv(13 downto 0);
      ptr_deref_941_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_gather_scatter
    process(type_cast_943_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_943_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_941_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_root_address_inst
    process(ptr_deref_941_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_941_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1312_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_880;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1312_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1312_branch_req_0,
          ack0 => if_stmt_1312_branch_ack_0,
          ack1 => if_stmt_1312_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1484_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1483;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1484_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1484_branch_req_0,
          ack0 => if_stmt_1484_branch_ack_0,
          ack1 => if_stmt_1484_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_421_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp513_420;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_421_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_421_branch_req_0,
          ack0 => if_stmt_421_branch_ack_0,
          ack1 => if_stmt_421_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_436_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194509_435;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_436_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_436_branch_req_0,
          ack0 => if_stmt_436_branch_ack_0,
          ack1 => if_stmt_436_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_637_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_636;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_637_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_637_branch_req_0,
          ack0 => if_stmt_637_branch_ack_0,
          ack1 => if_stmt_637_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_844_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_843;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_844_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_844_branch_req_0,
          ack0 => if_stmt_844_branch_ack_0,
          ack1 => if_stmt_844_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_881_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_880;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_881_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_881_branch_req_0,
          ack0 => if_stmt_881_branch_ack_0,
          ack1 => if_stmt_881_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_956_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_955;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_956_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_956_branch_req_0,
          ack0 => if_stmt_956_branch_ack_0,
          ack1 => if_stmt_956_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1335_inst
    process(tmp520_1324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp520_1324, type_cast_1334_wire_constant, tmp_var);
      tmp520x_xop_1336 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_257_inst
    process(add74_253, shr_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_253, shr_241, tmp_var);
      add79_258 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_453_inst
    process(shr_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_241, type_cast_452_wire_constant, tmp_var);
      tmp562x_xop_454 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_660_inst
    process(tmp548_649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp548_649, type_cast_659_wire_constant, tmp_var);
      tmp548x_xop_661 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_904_inst
    process(tmp532_893) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp532_893, type_cast_903_wire_constant, tmp_var);
      tmp532x_xop_905 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1345_inst
    process(iNsTr_196_1340) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_196_1340, type_cast_1344_wire_constant, tmp_var);
      xx_xop_1346 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1477_inst
    process(indvar_1356) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1356, type_cast_1476_wire_constant, tmp_var);
      indvarx_xnext_1478 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_463_inst
    process(iNsTr_26_458) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_458, type_cast_462_wire_constant, tmp_var);
      xx_xop571_464 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_630_inst
    process(indvar555_474) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar555_474, type_cast_629_wire_constant, tmp_var);
      indvarx_xnext556_631 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_670_inst
    process(iNsTr_39_665) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_665, type_cast_669_wire_constant, tmp_var);
      xx_xop570_671 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_837_inst
    process(indvar539_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar539_681, type_cast_836_wire_constant, tmp_var);
      indvarx_xnext540_838 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_914_inst
    process(iNsTr_53_909) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_909, type_cast_913_wire_constant, tmp_var);
      xx_xop569_915 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_949_inst
    process(indvar525_925) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar525_925, type_cast_948_wire_constant, tmp_var);
      indvarx_xnext526_950 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_252_inst
    process(iNsTr_14_247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_247, type_cast_251_wire_constant, tmp_var);
      add74_253 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1482_inst
    process(indvarx_xnext_1478, tmp524_1353) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1478, tmp524_1353, tmp_var);
      exitcond1_1483 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_635_inst
    process(indvarx_xnext556_631, tmp567_471) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext556_631, tmp567_471, tmp_var);
      exitcond3_636 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_842_inst
    process(indvarx_xnext540_838, tmp553_678) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext540_838, tmp553_678, tmp_var);
      exitcond2_843 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_954_inst
    process(indvarx_xnext526_950, tmp537_922) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext526_950, tmp537_922, tmp_var);
      exitcond_955 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1050_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_1049_wire_constant, tmp_var);
      shr304_1051 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1106_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_1105_wire_constant, tmp_var);
      shr321_1107 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1162_inst
    process(add79_258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_258, type_cast_1161_wire_constant, tmp_var);
      shr338_1163 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1323_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_874, type_cast_1322_wire_constant, tmp_var);
      tmp520_1324 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_240_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_239_wire_constant, tmp_var);
      shr_241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_246_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_245_wire_constant, tmp_var);
      iNsTr_14_247 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_648_inst
    process(mul91_289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_289, type_cast_647_wire_constant, tmp_var);
      tmp548_649 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_892_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_874, type_cast_891_wire_constant, tmp_var);
      tmp532_893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1221_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1220_wire_constant, tmp_var);
      shr364_1222 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1231_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1230_wire_constant, tmp_var);
      shr370_1232 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1241_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1240_wire_constant, tmp_var);
      shr376_1242 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1251_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1250_wire_constant, tmp_var);
      shr382_1252 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1261_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1260_wire_constant, tmp_var);
      shr388_1262 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1271_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1270_wire_constant, tmp_var);
      shr394_1272 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1281_inst
    process(sub_1212) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1212, type_cast_1280_wire_constant, tmp_var);
      shr400_1282 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1383_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1382_wire_constant, tmp_var);
      shr440_1384 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1393_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1392_wire_constant, tmp_var);
      shr446_1394 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1403_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1402_wire_constant, tmp_var);
      shr452_1404 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1413_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1412_wire_constant, tmp_var);
      shr458_1414 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1423_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1422_wire_constant, tmp_var);
      shr464_1424 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1433_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1432_wire_constant, tmp_var);
      shr470_1434 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1443_inst
    process(tmp433_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1374, type_cast_1442_wire_constant, tmp_var);
      shr476_1444 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(conv63_221, conv61_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_221, conv61_217, tmp_var);
      mul_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_234_inst
    process(mul_230, conv65_225) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_230, conv65_225, tmp_var);
      mul66_235 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_278_inst
    process(conv84_266, conv82_262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_266, conv82_262, tmp_var);
      mul85_279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_283_inst
    process(mul85_279, conv87_270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_279, conv87_270, tmp_var);
      mul88_284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_288_inst
    process(mul88_284, conv90_274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_284, conv90_274, tmp_var);
      mul91_289 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_868_inst
    process(conv255_860, conv253_856) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_860, conv253_856, tmp_var);
      mul256_869 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_873_inst
    process(mul256_869, conv258_864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_869, conv258_864, tmp_var);
      mul259_874 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_112_inst
    process(shl18_101, conv20_108) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_101, conv20_108, tmp_var);
      add21_113 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_137_inst
    process(shl27_126, conv29_133) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_126, conv29_133, tmp_var);
      add30_138 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_162_inst
    process(shl36_151, conv38_158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_151, conv38_158, tmp_var);
      add39_163 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_187_inst
    process(shl45_176, conv47_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_176, conv47_183, tmp_var);
      add48_188 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_212_inst
    process(shl54_201, conv56_208) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_201, conv56_208, tmp_var);
      add57_213 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_313_inst
    process(shl96_302, conv98_309) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_302, conv98_309, tmp_var);
      add99_314 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_338_inst
    process(shl105_327, conv107_334) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_327, conv107_334, tmp_var);
      add108_339 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_363_inst
    process(shl114_352, conv116_359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_352, conv116_359, tmp_var);
      add117_364 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_388_inst
    process(shl123_377, conv125_384) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_377, conv125_384, tmp_var);
      add126_389 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_413_inst
    process(shl132_402, conv134_409) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_402, conv134_409, tmp_var);
      add135_414 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_62_inst
    process(shl_51, conv3_58) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_51, conv3_58, tmp_var);
      add_63 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_87_inst
    process(shl9_76, conv11_83) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_76, conv11_83, tmp_var);
      add12_88 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_512_inst
    process(shl146_501, conv149_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_501, conv149_508, tmp_var);
      add150_513 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_530_inst
    process(shl152_519, conv155_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_519, conv155_526, tmp_var);
      add156_531 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_548_inst
    process(shl158_537, conv161_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_537, conv161_544, tmp_var);
      add162_549 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_566_inst
    process(shl164_555, conv167_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_555, conv167_562, tmp_var);
      add168_567 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_584_inst
    process(shl170_573, conv173_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_573, conv173_580, tmp_var);
      add174_585 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_602_inst
    process(shl176_591, conv179_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_591, conv179_598, tmp_var);
      add180_603 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_620_inst
    process(shl182_609, conv185_616) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_609, conv185_616, tmp_var);
      add186_621 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_719_inst
    process(shl202_708, conv205_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_708, conv205_715, tmp_var);
      add206_720 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_737_inst
    process(shl208_726, conv211_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_726, conv211_733, tmp_var);
      add212_738 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_755_inst
    process(shl214_744, conv217_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_744, conv217_751, tmp_var);
      add218_756 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_773_inst
    process(shl220_762, conv223_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_762, conv223_769, tmp_var);
      add224_774 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_791_inst
    process(shl226_780, conv229_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_780, conv229_787, tmp_var);
      add230_792 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_809_inst
    process(shl232_798, conv235_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_798, conv235_805, tmp_var);
      add236_810 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_827_inst
    process(shl238_816, conv241_823) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_816, conv241_823, tmp_var);
      add242_828 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_100_inst
    process(conv17_95) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_95, type_cast_99_wire_constant, tmp_var);
      shl18_101 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_125_inst
    process(conv26_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_120, type_cast_124_wire_constant, tmp_var);
      shl27_126 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_150_inst
    process(conv35_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_145, type_cast_149_wire_constant, tmp_var);
      shl36_151 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_175_inst
    process(conv44_170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_170, type_cast_174_wire_constant, tmp_var);
      shl45_176 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_200_inst
    process(conv53_195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_195, type_cast_199_wire_constant, tmp_var);
      shl54_201 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_301_inst
    process(conv95_296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_296, type_cast_300_wire_constant, tmp_var);
      shl96_302 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_326_inst
    process(conv104_321) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_321, type_cast_325_wire_constant, tmp_var);
      shl105_327 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_351_inst
    process(conv113_346) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_346, type_cast_350_wire_constant, tmp_var);
      shl114_352 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_376_inst
    process(conv122_371) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_371, type_cast_375_wire_constant, tmp_var);
      shl123_377 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_401_inst
    process(conv131_396) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_396, type_cast_400_wire_constant, tmp_var);
      shl132_402 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_50_inst
    process(conv1_45) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_45, type_cast_49_wire_constant, tmp_var);
      shl_51 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_75_inst
    process(conv8_70) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_70, type_cast_74_wire_constant, tmp_var);
      shl9_76 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_500_inst
    process(conv144_495) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_495, type_cast_499_wire_constant, tmp_var);
      shl146_501 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_518_inst
    process(add150_513) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_513, type_cast_517_wire_constant, tmp_var);
      shl152_519 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_536_inst
    process(add156_531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_531, type_cast_535_wire_constant, tmp_var);
      shl158_537 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_554_inst
    process(add162_549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_549, type_cast_553_wire_constant, tmp_var);
      shl164_555 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_572_inst
    process(add168_567) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_567, type_cast_571_wire_constant, tmp_var);
      shl170_573 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_590_inst
    process(add174_585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_585, type_cast_589_wire_constant, tmp_var);
      shl176_591 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_608_inst
    process(add180_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_603, type_cast_607_wire_constant, tmp_var);
      shl182_609 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_707_inst
    process(conv200_702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_702, type_cast_706_wire_constant, tmp_var);
      shl202_708 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_725_inst
    process(add206_720) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_720, type_cast_724_wire_constant, tmp_var);
      shl208_726 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_743_inst
    process(add212_738) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_738, type_cast_742_wire_constant, tmp_var);
      shl214_744 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_761_inst
    process(add218_756) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_756, type_cast_760_wire_constant, tmp_var);
      shl220_762 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_779_inst
    process(add224_774) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_774, type_cast_778_wire_constant, tmp_var);
      shl226_780 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_797_inst
    process(add230_792) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_792, type_cast_796_wire_constant, tmp_var);
      shl232_798 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_815_inst
    process(add236_810) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_810, type_cast_814_wire_constant, tmp_var);
      shl238_816 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1211_inst
    process(conv355_1207, conv276_973) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1207, conv276_973, tmp_var);
      sub_1212 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1329_inst
    process(tmp520_1324) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp520_1324, type_cast_1328_wire_constant, tmp_var);
      tmp521_1330 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_419_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_235, type_cast_418_wire_constant, tmp_var);
      cmp513_420 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_434_inst
    process(mul91_289) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_289, type_cast_433_wire_constant, tmp_var);
      cmp194509_435 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_447_inst
    process(shr_241) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_241, type_cast_446_wire_constant, tmp_var);
      tmp563_448 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_654_inst
    process(tmp548_649) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp548_649, type_cast_653_wire_constant, tmp_var);
      tmp549_655 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_879_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_874, type_cast_878_wire_constant, tmp_var);
      cmp264505_880 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_898_inst
    process(tmp532_893) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp532_893, type_cast_897_wire_constant, tmp_var);
      tmp533_899 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1368_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1367_scaled;
      array_obj_ref_1368_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1368_index_offset_req_0;
      array_obj_ref_1368_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1368_index_offset_req_1;
      array_obj_ref_1368_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_486_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar555_485_scaled;
      array_obj_ref_486_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_486_index_offset_req_0;
      array_obj_ref_486_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_486_index_offset_req_1;
      array_obj_ref_486_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_693_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar539_692_scaled;
      array_obj_ref_693_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_693_index_offset_req_0;
      array_obj_ref_693_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_693_index_offset_req_1;
      array_obj_ref_693_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_937_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar525_936_scaled;
      array_obj_ref_937_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_937_index_offset_req_0;
      array_obj_ref_937_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_937_index_offset_req_1;
      array_obj_ref_937_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1205_inst
    process(call354_1202) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1202, tmp_var);
      type_cast_1205_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_971_inst
    process(call275_967) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_967, tmp_var);
      type_cast_971_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1373_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1373_load_0_req_0;
      ptr_deref_1373_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1373_load_0_req_1;
      ptr_deref_1373_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1373_word_address_0;
      ptr_deref_1373_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_623_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_623_store_0_req_0;
      ptr_deref_623_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_623_store_0_req_1;
      ptr_deref_623_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_623_word_address_0;
      data_in <= ptr_deref_623_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_830_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_830_store_0_req_0;
      ptr_deref_830_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_830_store_0_req_1;
      ptr_deref_830_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_830_word_address_0;
      data_in <= ptr_deref_830_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(10 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_941_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_941_store_0_req_0;
      ptr_deref_941_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_941_store_0_req_1;
      ptr_deref_941_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_941_word_address_0;
      data_in <= ptr_deref_941_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1189_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1189_inst_req_0;
      RPIPE_Block0_done_1189_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1189_inst_req_1;
      RPIPE_Block0_done_1189_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1190 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1192_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1192_inst_req_0;
      RPIPE_Block1_done_1192_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1192_inst_req_1;
      RPIPE_Block1_done_1192_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1193 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1195_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1195_inst_req_0;
      RPIPE_Block2_done_1195_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1195_inst_req_1;
      RPIPE_Block2_done_1195_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1196 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1198_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1198_inst_req_0;
      RPIPE_Block3_done_1198_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1198_inst_req_1;
      RPIPE_Block3_done_1198_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1199 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_53_inst RPIPE_ConvTranspose_input_pipe_40_inst RPIPE_ConvTranspose_input_pipe_710_inst RPIPE_ConvTranspose_input_pipe_128_inst RPIPE_ConvTranspose_input_pipe_697_inst RPIPE_ConvTranspose_input_pipe_818_inst RPIPE_ConvTranspose_input_pipe_782_inst RPIPE_ConvTranspose_input_pipe_728_inst RPIPE_ConvTranspose_input_pipe_153_inst RPIPE_ConvTranspose_input_pipe_178_inst RPIPE_ConvTranspose_input_pipe_140_inst RPIPE_ConvTranspose_input_pipe_800_inst RPIPE_ConvTranspose_input_pipe_115_inst RPIPE_ConvTranspose_input_pipe_78_inst RPIPE_ConvTranspose_input_pipe_746_inst RPIPE_ConvTranspose_input_pipe_165_inst RPIPE_ConvTranspose_input_pipe_764_inst RPIPE_ConvTranspose_input_pipe_90_inst RPIPE_ConvTranspose_input_pipe_103_inst RPIPE_ConvTranspose_input_pipe_65_inst RPIPE_ConvTranspose_input_pipe_190_inst RPIPE_ConvTranspose_input_pipe_203_inst RPIPE_ConvTranspose_input_pipe_291_inst RPIPE_ConvTranspose_input_pipe_304_inst RPIPE_ConvTranspose_input_pipe_316_inst RPIPE_ConvTranspose_input_pipe_329_inst RPIPE_ConvTranspose_input_pipe_341_inst RPIPE_ConvTranspose_input_pipe_354_inst RPIPE_ConvTranspose_input_pipe_366_inst RPIPE_ConvTranspose_input_pipe_379_inst RPIPE_ConvTranspose_input_pipe_391_inst RPIPE_ConvTranspose_input_pipe_404_inst RPIPE_ConvTranspose_input_pipe_490_inst RPIPE_ConvTranspose_input_pipe_503_inst RPIPE_ConvTranspose_input_pipe_521_inst RPIPE_ConvTranspose_input_pipe_539_inst RPIPE_ConvTranspose_input_pipe_557_inst RPIPE_ConvTranspose_input_pipe_575_inst RPIPE_ConvTranspose_input_pipe_593_inst RPIPE_ConvTranspose_input_pipe_611_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_710_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_697_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_818_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_782_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_800_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_746_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_764_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_304_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_379_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_404_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_490_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_503_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_521_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_539_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_575_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_710_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_697_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_818_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_782_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_800_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_746_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_764_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_304_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_379_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_404_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_490_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_503_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_521_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_539_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_575_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_710_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_697_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_818_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_782_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_800_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_746_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_764_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_304_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_379_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_404_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_490_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_503_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_521_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_539_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_575_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_710_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_697_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_818_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_782_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_800_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_746_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_764_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_304_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_379_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_404_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_490_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_503_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_521_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_539_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_575_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call2_54 <= data_out(319 downto 312);
      call_41 <= data_out(311 downto 304);
      call203_711 <= data_out(303 downto 296);
      call28_129 <= data_out(295 downto 288);
      call199_698 <= data_out(287 downto 280);
      call239_819 <= data_out(279 downto 272);
      call227_783 <= data_out(271 downto 264);
      call209_729 <= data_out(263 downto 256);
      call37_154 <= data_out(255 downto 248);
      call46_179 <= data_out(247 downto 240);
      call32_141 <= data_out(239 downto 232);
      call233_801 <= data_out(231 downto 224);
      call23_116 <= data_out(223 downto 216);
      call10_79 <= data_out(215 downto 208);
      call215_747 <= data_out(207 downto 200);
      call41_166 <= data_out(199 downto 192);
      call221_765 <= data_out(191 downto 184);
      call14_91 <= data_out(183 downto 176);
      call19_104 <= data_out(175 downto 168);
      call5_66 <= data_out(167 downto 160);
      call50_191 <= data_out(159 downto 152);
      call55_204 <= data_out(151 downto 144);
      call92_292 <= data_out(143 downto 136);
      call97_305 <= data_out(135 downto 128);
      call101_317 <= data_out(127 downto 120);
      call106_330 <= data_out(119 downto 112);
      call110_342 <= data_out(111 downto 104);
      call115_355 <= data_out(103 downto 96);
      call119_367 <= data_out(95 downto 88);
      call124_380 <= data_out(87 downto 80);
      call128_392 <= data_out(79 downto 72);
      call133_405 <= data_out(71 downto 64);
      call143_491 <= data_out(63 downto 56);
      call147_504 <= data_out(55 downto 48);
      call153_522 <= data_out(47 downto 40);
      call159_540 <= data_out(39 downto 32);
      call165_558 <= data_out(31 downto 24);
      call171_576 <= data_out(23 downto 16);
      call177_594 <= data_out(15 downto 8);
      call183_612 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_1013_inst WPIPE_Block0_start_975_inst WPIPE_Block0_start_978_inst WPIPE_Block0_start_981_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_993_inst WPIPE_Block0_start_996_inst WPIPE_Block0_start_999_inst WPIPE_Block0_start_984_inst WPIPE_Block0_start_1002_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_1006_inst WPIPE_Block0_start_1010_inst WPIPE_Block0_start_1016_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_1013_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_975_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_981_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_993_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_996_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_999_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_984_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_1002_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_1006_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_1010_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_1016_inst_req_0;
      WPIPE_Block0_start_1013_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_975_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_981_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_993_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_996_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_999_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_984_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_1002_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_1006_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_1010_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_1016_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_1013_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_975_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_981_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_993_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_996_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_999_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_984_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_1002_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_1006_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_1010_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_1016_inst_req_1;
      WPIPE_Block0_start_1013_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_975_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_981_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_993_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_996_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_999_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_984_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_1002_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_1006_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_1010_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_1016_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add126_389 & add_63 & add12_88 & add21_113 & add48_188 & add57_213 & add99_314 & add108_339 & add30_138 & type_cast_1004_wire_constant & add39_163 & type_cast_1008_wire_constant & add117_364 & add135_414;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1056_inst WPIPE_Block1_start_1022_inst WPIPE_Block1_start_1063_inst WPIPE_Block1_start_1066_inst WPIPE_Block1_start_1031_inst WPIPE_Block1_start_1034_inst WPIPE_Block1_start_1069_inst WPIPE_Block1_start_1025_inst WPIPE_Block1_start_1072_inst WPIPE_Block1_start_1037_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1028_inst WPIPE_Block1_start_1040_inst WPIPE_Block1_start_1043_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1056_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1022_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1063_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1031_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1034_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1069_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1025_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1072_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1037_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1028_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1040_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1043_inst_req_0;
      WPIPE_Block1_start_1056_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1063_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1031_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1034_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1069_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1025_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1072_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1037_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1028_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1040_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1043_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1056_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1022_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1063_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1031_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1034_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1069_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1025_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1072_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1037_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1028_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1040_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1043_inst_req_1;
      WPIPE_Block1_start_1056_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1063_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1031_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1034_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1069_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1025_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1072_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1037_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1028_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1040_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1043_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv305_1055 & add12_88 & conv307_1062 & add117_364 & add39_163 & add48_188 & add126_389 & add21_113 & add135_414 & add57_213 & add_63 & add30_138 & add99_314 & add108_339;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1090_inst WPIPE_Block2_start_1112_inst WPIPE_Block2_start_1128_inst WPIPE_Block2_start_1087_inst WPIPE_Block2_start_1093_inst WPIPE_Block2_start_1096_inst WPIPE_Block2_start_1084_inst WPIPE_Block2_start_1099_inst WPIPE_Block2_start_1075_inst WPIPE_Block2_start_1078_inst WPIPE_Block2_start_1081_inst WPIPE_Block2_start_1119_inst WPIPE_Block2_start_1122_inst WPIPE_Block2_start_1125_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1090_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1112_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1128_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1087_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1093_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1096_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1084_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1099_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1075_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1078_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1081_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1119_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1122_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1125_inst_req_0;
      WPIPE_Block2_start_1090_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1112_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1128_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1087_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1093_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1096_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1084_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1099_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1075_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1078_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1081_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1119_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1122_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1125_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1090_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1112_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1128_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1087_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1093_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1096_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1084_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1099_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1075_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1078_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1081_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1119_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1122_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1125_inst_req_1;
      WPIPE_Block2_start_1090_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1112_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1128_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1087_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1093_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1096_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1084_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1099_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1075_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1078_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1081_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1119_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1122_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1125_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add48_188 & conv322_1111 & add135_414 & add39_163 & add57_213 & add99_314 & add30_138 & add108_339 & add_63 & add12_88 & add21_113 & conv324_1118 & add117_364 & add126_389;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1134_inst WPIPE_Block3_start_1149_inst WPIPE_Block3_start_1178_inst WPIPE_Block3_start_1131_inst WPIPE_Block3_start_1137_inst WPIPE_Block3_start_1143_inst WPIPE_Block3_start_1152_inst WPIPE_Block3_start_1140_inst WPIPE_Block3_start_1168_inst WPIPE_Block3_start_1181_inst WPIPE_Block3_start_1155_inst WPIPE_Block3_start_1146_inst WPIPE_Block3_start_1184_inst WPIPE_Block3_start_1175_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1134_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1149_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1178_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1131_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1137_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1143_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1152_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1140_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1168_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1181_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1155_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1146_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1184_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1175_inst_req_0;
      WPIPE_Block3_start_1134_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1149_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1178_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1131_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1137_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1143_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1152_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1140_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1168_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1181_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1155_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1146_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1184_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1175_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1134_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1149_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1178_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1131_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1137_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1143_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1152_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1140_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1168_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1181_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1155_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1146_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1184_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1175_inst_req_1;
      WPIPE_Block3_start_1134_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1149_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1178_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1131_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1137_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1143_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1152_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1140_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1168_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1181_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1155_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1146_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1184_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1175_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add12_88 & add57_213 & add117_364 & add_63 & add21_113 & add39_163 & add99_314 & add30_138 & conv339_1167 & add126_389 & add108_339 & add48_188 & add135_414 & conv341_1174;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1302_inst WPIPE_ConvTranspose_output_pipe_1299_inst WPIPE_ConvTranspose_output_pipe_1296_inst WPIPE_ConvTranspose_output_pipe_1287_inst WPIPE_ConvTranspose_output_pipe_1293_inst WPIPE_ConvTranspose_output_pipe_1290_inst WPIPE_ConvTranspose_output_pipe_1308_inst WPIPE_ConvTranspose_output_pipe_1305_inst WPIPE_ConvTranspose_output_pipe_1449_inst WPIPE_ConvTranspose_output_pipe_1452_inst WPIPE_ConvTranspose_output_pipe_1455_inst WPIPE_ConvTranspose_output_pipe_1458_inst WPIPE_ConvTranspose_output_pipe_1461_inst WPIPE_ConvTranspose_output_pipe_1464_inst WPIPE_ConvTranspose_output_pipe_1467_inst WPIPE_ConvTranspose_output_pipe_1470_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1308_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1305_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1449_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1452_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1455_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1458_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1461_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1464_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1467_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1470_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1308_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1305_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1449_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1452_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1455_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1458_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1461_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1464_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1467_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1470_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1302_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1299_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1296_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1287_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1293_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1290_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1308_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1305_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1449_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1452_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1455_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1458_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1461_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1464_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1467_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1470_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1302_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1299_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1296_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1287_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1293_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1290_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1308_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1305_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1449_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1452_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1455_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1458_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1461_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1464_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1467_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1470_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv373_1236 & conv379_1246 & conv385_1256 & conv403_1286 & conv391_1266 & conv397_1276 & conv361_1216 & conv367_1226 & conv479_1448 & conv473_1438 & conv467_1428 & conv461_1418 & conv455_1408 & conv449_1398 & conv443_1388 & conv437_1378;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1202_call call_stmt_967_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1202_call_req_0;
      reqL_unguarded(0) <= call_stmt_967_call_req_0;
      call_stmt_1202_call_ack_0 <= ackL_unguarded(1);
      call_stmt_967_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1202_call_req_1;
      reqR_unguarded(0) <= call_stmt_967_call_req_1;
      call_stmt_1202_call_ack_1 <= ackR_unguarded(1);
      call_stmt_967_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call354_1202 <= data_out(127 downto 64);
      call275_967 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3763_start: Boolean;
  signal convTransposeA_CP_3763_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1512_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_ack_0 : boolean;
  signal type_cast_1789_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1500_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1524_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1500_inst_req_1 : boolean;
  signal W_input_dim1x_x1_1790_delayed_2_0_1797_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1503_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1500_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1524_inst_req_0 : boolean;
  signal addr_of_1748_final_reg_ack_0 : boolean;
  signal W_input_dim1x_x1_1790_delayed_2_0_1797_inst_ack_0 : boolean;
  signal ptr_deref_1754_store_0_ack_1 : boolean;
  signal RPIPE_Block0_start_1524_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1540_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1558_inst_req_1 : boolean;
  signal W_add96_1773_delayed_1_0_1777_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1558_inst_ack_1 : boolean;
  signal ptr_deref_1729_load_0_ack_1 : boolean;
  signal type_cast_1759_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1512_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1503_inst_req_1 : boolean;
  signal array_obj_ref_1747_index_offset_ack_1 : boolean;
  signal RPIPE_Block0_start_1558_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1540_inst_ack_0 : boolean;
  signal type_cast_1789_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1555_inst_req_0 : boolean;
  signal W_add96_1773_delayed_1_0_1777_inst_ack_1 : boolean;
  signal type_cast_1531_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_1 : boolean;
  signal ptr_deref_1729_load_0_req_1 : boolean;
  signal array_obj_ref_1747_index_offset_req_0 : boolean;
  signal type_cast_1531_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_0 : boolean;
  signal array_obj_ref_1747_index_offset_ack_0 : boolean;
  signal RPIPE_Block0_start_1555_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1558_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1540_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1540_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1506_inst_req_1 : boolean;
  signal type_cast_1544_inst_ack_1 : boolean;
  signal type_cast_1763_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1512_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1521_inst_req_0 : boolean;
  signal type_cast_1763_inst_req_1 : boolean;
  signal addr_of_1748_final_reg_req_0 : boolean;
  signal do_while_stmt_1636_branch_ack_1 : boolean;
  signal RPIPE_Block0_start_1555_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1524_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1506_inst_req_0 : boolean;
  signal type_cast_1759_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1518_inst_req_0 : boolean;
  signal type_cast_1759_inst_req_0 : boolean;
  signal type_cast_1544_inst_req_0 : boolean;
  signal if_stmt_1850_branch_ack_0 : boolean;
  signal RPIPE_Block0_start_1503_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1506_inst_ack_0 : boolean;
  signal type_cast_1544_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1512_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1518_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1503_inst_ack_0 : boolean;
  signal type_cast_1531_inst_req_1 : boolean;
  signal type_cast_1531_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1515_inst_ack_1 : boolean;
  signal type_cast_1763_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1555_inst_ack_0 : boolean;
  signal addr_of_1748_final_reg_req_1 : boolean;
  signal if_stmt_1850_branch_ack_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1521_inst_ack_1 : boolean;
  signal addr_of_1748_final_reg_ack_1 : boolean;
  signal type_cast_1544_inst_req_1 : boolean;
  signal ptr_deref_1754_store_0_req_1 : boolean;
  signal type_cast_1759_inst_req_1 : boolean;
  signal type_cast_1763_inst_ack_0 : boolean;
  signal type_cast_1601_inst_req_1 : boolean;
  signal W_add96_1773_delayed_1_0_1777_inst_req_0 : boolean;
  signal type_cast_1601_inst_ack_1 : boolean;
  signal type_cast_1601_inst_req_0 : boolean;
  signal W_add96_1773_delayed_1_0_1777_inst_ack_0 : boolean;
  signal type_cast_1601_inst_ack_0 : boolean;
  signal if_stmt_1850_branch_req_0 : boolean;
  signal array_obj_ref_1747_index_offset_req_1 : boolean;
  signal type_cast_1585_inst_req_0 : boolean;
  signal type_cast_1589_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1552_inst_ack_1 : boolean;
  signal W_input_dim0x_x1_1804_delayed_3_0_1814_inst_req_1 : boolean;
  signal type_cast_1589_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1552_inst_req_1 : boolean;
  signal W_input_dim1x_x1_1790_delayed_2_0_1797_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1527_inst_ack_1 : boolean;
  signal type_cast_1589_inst_req_0 : boolean;
  signal type_cast_1589_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1527_inst_req_1 : boolean;
  signal ptr_deref_1754_store_0_ack_0 : boolean;
  signal ptr_deref_1754_store_0_req_0 : boolean;
  signal RPIPE_Block0_start_1552_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1552_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1527_inst_ack_0 : boolean;
  signal W_input_dim0x_x1_1804_delayed_3_0_1814_inst_ack_1 : boolean;
  signal type_cast_1585_inst_req_1 : boolean;
  signal type_cast_1585_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1527_inst_req_0 : boolean;
  signal type_cast_1585_inst_ack_0 : boolean;
  signal type_cast_1605_inst_req_0 : boolean;
  signal type_cast_1605_inst_ack_0 : boolean;
  signal type_cast_1605_inst_req_1 : boolean;
  signal type_cast_1605_inst_ack_1 : boolean;
  signal ptr_deref_1729_load_0_ack_0 : boolean;
  signal do_while_stmt_1636_branch_req_0 : boolean;
  signal type_cast_1812_inst_ack_1 : boolean;
  signal type_cast_1812_inst_req_1 : boolean;
  signal W_input_dim1x_x1_1790_delayed_2_0_1797_inst_ack_1 : boolean;
  signal do_while_stmt_1636_branch_ack_0 : boolean;
  signal type_cast_1789_inst_ack_1 : boolean;
  signal phi_stmt_1638_req_0 : boolean;
  signal type_cast_1831_inst_ack_1 : boolean;
  signal type_cast_1831_inst_req_1 : boolean;
  signal phi_stmt_1638_req_1 : boolean;
  signal type_cast_1812_inst_ack_0 : boolean;
  signal phi_stmt_1638_ack_0 : boolean;
  signal type_cast_1831_inst_ack_0 : boolean;
  signal W_input_dim0x_x1_1804_delayed_3_0_1814_inst_ack_0 : boolean;
  signal type_cast_1641_inst_req_0 : boolean;
  signal type_cast_1641_inst_ack_0 : boolean;
  signal ptr_deref_1729_load_0_req_0 : boolean;
  signal W_input_dim0x_x1_1804_delayed_3_0_1814_inst_req_0 : boolean;
  signal type_cast_1641_inst_req_1 : boolean;
  signal type_cast_1641_inst_ack_1 : boolean;
  signal type_cast_1789_inst_req_1 : boolean;
  signal type_cast_1812_inst_req_0 : boolean;
  signal W_arrayidx81_1750_delayed_6_0_1750_inst_ack_1 : boolean;
  signal W_arrayidx81_1750_delayed_6_0_1750_inst_req_1 : boolean;
  signal type_cast_1831_inst_req_0 : boolean;
  signal W_arrayidx81_1750_delayed_6_0_1750_inst_ack_0 : boolean;
  signal W_arrayidx81_1750_delayed_6_0_1750_inst_req_0 : boolean;
  signal phi_stmt_1643_req_0 : boolean;
  signal phi_stmt_1643_req_1 : boolean;
  signal phi_stmt_1643_ack_0 : boolean;
  signal type_cast_1646_inst_req_0 : boolean;
  signal type_cast_1646_inst_ack_0 : boolean;
  signal type_cast_1646_inst_req_1 : boolean;
  signal type_cast_1646_inst_ack_1 : boolean;
  signal phi_stmt_1648_req_0 : boolean;
  signal phi_stmt_1648_req_1 : boolean;
  signal phi_stmt_1648_ack_0 : boolean;
  signal type_cast_1651_inst_req_0 : boolean;
  signal type_cast_1651_inst_ack_0 : boolean;
  signal type_cast_1651_inst_req_1 : boolean;
  signal type_cast_1651_inst_ack_1 : boolean;
  signal phi_stmt_1653_req_0 : boolean;
  signal phi_stmt_1653_req_1 : boolean;
  signal phi_stmt_1653_ack_0 : boolean;
  signal type_cast_1656_inst_req_0 : boolean;
  signal type_cast_1656_inst_ack_0 : boolean;
  signal type_cast_1656_inst_req_1 : boolean;
  signal type_cast_1656_inst_ack_1 : boolean;
  signal type_cast_1686_inst_req_0 : boolean;
  signal type_cast_1686_inst_ack_0 : boolean;
  signal type_cast_1686_inst_req_1 : boolean;
  signal type_cast_1686_inst_ack_1 : boolean;
  signal type_cast_1690_inst_req_0 : boolean;
  signal type_cast_1690_inst_ack_0 : boolean;
  signal type_cast_1690_inst_req_1 : boolean;
  signal type_cast_1690_inst_ack_1 : boolean;
  signal type_cast_1694_inst_req_0 : boolean;
  signal type_cast_1694_inst_ack_0 : boolean;
  signal type_cast_1694_inst_req_1 : boolean;
  signal type_cast_1694_inst_ack_1 : boolean;
  signal type_cast_1718_inst_req_0 : boolean;
  signal type_cast_1718_inst_ack_0 : boolean;
  signal type_cast_1718_inst_req_1 : boolean;
  signal type_cast_1718_inst_ack_1 : boolean;
  signal array_obj_ref_1724_index_offset_req_0 : boolean;
  signal array_obj_ref_1724_index_offset_ack_0 : boolean;
  signal array_obj_ref_1724_index_offset_req_1 : boolean;
  signal array_obj_ref_1724_index_offset_ack_1 : boolean;
  signal addr_of_1725_final_reg_req_0 : boolean;
  signal addr_of_1725_final_reg_ack_0 : boolean;
  signal addr_of_1725_final_reg_req_1 : boolean;
  signal addr_of_1725_final_reg_ack_1 : boolean;
  signal WPIPE_Block0_done_1856_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1856_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1856_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1856_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3763_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3763_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3763: Block -- control-path 
    signal convTransposeA_CP_3763_elements: BooleanArray(222 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3763_elements(0) <= convTransposeA_CP_3763_start;
    convTransposeA_CP_3763_symbol <= convTransposeA_CP_3763_elements(222);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559__entry__
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/branch_block_stmt_1498__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/cr
      -- 
    rr_3797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => RPIPE_Block0_start_1500_inst_req_0); -- 
    cr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => type_cast_1531_inst_req_1); -- 
    cr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(0), ack => type_cast_1544_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	218 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	219 
    -- CP-element group 1: 	220 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850__entry__
      -- CP-element group 1: 	 branch_block_stmt_1498/do_while_stmt_1636__exit__
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/if_stmt_1850_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1498/R_whilex_xbody_whilex_xend_taken_1851_place
      -- 
    branch_req_4660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(1), ack => if_stmt_1850_branch_req_0); -- 
    convTransposeA_CP_3763_elements(1) <= convTransposeA_CP_3763_elements(218);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_update_start_
      -- 
    ra_3798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1500_inst_ack_0, ack => convTransposeA_CP_3763_elements(2)); -- 
    cr_3802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(2), ack => RPIPE_Block0_start_1500_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1500_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/rr
      -- 
    ca_3803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1500_inst_ack_1, ack => convTransposeA_CP_3763_elements(3)); -- 
    rr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(3), ack => RPIPE_Block0_start_1503_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/$entry
      -- 
    ra_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1503_inst_ack_0, ack => convTransposeA_CP_3763_elements(4)); -- 
    cr_3816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(4), ack => RPIPE_Block0_start_1503_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1503_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_sample_start_
      -- 
    ca_3817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1503_inst_ack_1, ack => convTransposeA_CP_3763_elements(5)); -- 
    rr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(5), ack => RPIPE_Block0_start_1506_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Sample/ra
      -- 
    ra_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1506_inst_ack_0, ack => convTransposeA_CP_3763_elements(6)); -- 
    cr_3830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(6), ack => RPIPE_Block0_start_1506_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1506_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/rr
      -- 
    ca_3831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1506_inst_ack_1, ack => convTransposeA_CP_3763_elements(7)); -- 
    rr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(7), ack => RPIPE_Block0_start_1509_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/$entry
      -- 
    ra_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_0, ack => convTransposeA_CP_3763_elements(8)); -- 
    cr_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(8), ack => RPIPE_Block0_start_1509_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1509_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/$entry
      -- 
    ca_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_1, ack => convTransposeA_CP_3763_elements(9)); -- 
    rr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(9), ack => RPIPE_Block0_start_1512_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_update_start_
      -- 
    ra_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1512_inst_ack_0, ack => convTransposeA_CP_3763_elements(10)); -- 
    cr_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(10), ack => RPIPE_Block0_start_1512_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1512_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/$entry
      -- 
    ca_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1512_inst_ack_1, ack => convTransposeA_CP_3763_elements(11)); -- 
    rr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(11), ack => RPIPE_Block0_start_1515_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Sample/$exit
      -- 
    ra_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1515_inst_ack_0, ack => convTransposeA_CP_3763_elements(12)); -- 
    cr_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(12), ack => RPIPE_Block0_start_1515_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1515_Update/ca
      -- 
    ca_3873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1515_inst_ack_1, ack => convTransposeA_CP_3763_elements(13)); -- 
    rr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(13), ack => RPIPE_Block0_start_1518_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/$entry
      -- 
    ra_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1518_inst_ack_0, ack => convTransposeA_CP_3763_elements(14)); -- 
    cr_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(14), ack => RPIPE_Block0_start_1518_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1518_Update/$exit
      -- 
    ca_3887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1518_inst_ack_1, ack => convTransposeA_CP_3763_elements(15)); -- 
    rr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(15), ack => RPIPE_Block0_start_1521_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/cr
      -- 
    ra_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1521_inst_ack_0, ack => convTransposeA_CP_3763_elements(16)); -- 
    cr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(16), ack => RPIPE_Block0_start_1521_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1521_Update/ca
      -- 
    ca_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1521_inst_ack_1, ack => convTransposeA_CP_3763_elements(17)); -- 
    rr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(17), ack => RPIPE_Block0_start_1524_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Sample/ra
      -- 
    ra_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1524_inst_ack_0, ack => convTransposeA_CP_3763_elements(18)); -- 
    cr_3914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(18), ack => RPIPE_Block0_start_1524_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1524_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/$entry
      -- 
    ca_3915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1524_inst_ack_1, ack => convTransposeA_CP_3763_elements(19)); -- 
    rr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(19), ack => RPIPE_Block0_start_1527_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Sample/$exit
      -- 
    ra_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1527_inst_ack_0, ack => convTransposeA_CP_3763_elements(20)); -- 
    cr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(20), ack => RPIPE_Block0_start_1527_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1527_Update/$exit
      -- 
    ca_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1527_inst_ack_1, ack => convTransposeA_CP_3763_elements(21)); -- 
    rr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(21), ack => type_cast_1531_inst_req_0); -- 
    rr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(21), ack => RPIPE_Block0_start_1540_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_sample_completed_
      -- 
    ra_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_0, ack => convTransposeA_CP_3763_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1531_Update/ca
      -- 
    ca_3943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1531_inst_ack_1, ack => convTransposeA_CP_3763_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/$entry
      -- 
    ra_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1540_inst_ack_0, ack => convTransposeA_CP_3763_elements(24)); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(24), ack => RPIPE_Block0_start_1540_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1540_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/$entry
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1540_inst_ack_1, ack => convTransposeA_CP_3763_elements(25)); -- 
    rr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(25), ack => type_cast_1544_inst_req_0); -- 
    rr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(25), ack => RPIPE_Block0_start_1552_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Sample/ra
      -- 
    ra_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_0, ack => convTransposeA_CP_3763_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/type_cast_1544_Update/$exit
      -- 
    ca_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_1, ack => convTransposeA_CP_3763_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Sample/$exit
      -- 
    ra_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1552_inst_ack_0, ack => convTransposeA_CP_3763_elements(28)); -- 
    cr_3984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(28), ack => RPIPE_Block0_start_1552_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1552_update_completed_
      -- 
    ca_3985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1552_inst_ack_1, ack => convTransposeA_CP_3763_elements(29)); -- 
    rr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(29), ack => RPIPE_Block0_start_1555_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_sample_completed_
      -- 
    ra_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1555_inst_ack_0, ack => convTransposeA_CP_3763_elements(30)); -- 
    cr_3998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(30), ack => RPIPE_Block0_start_1555_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1555_update_completed_
      -- 
    ca_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1555_inst_ack_1, ack => convTransposeA_CP_3763_elements(31)); -- 
    rr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(31), ack => RPIPE_Block0_start_1558_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_sample_completed_
      -- 
    ra_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1558_inst_ack_0, ack => convTransposeA_CP_3763_elements(32)); -- 
    cr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(32), ack => RPIPE_Block0_start_1558_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/RPIPE_Block0_start_1558_Update/$exit
      -- 
    ca_4013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1558_inst_ack_1, ack => convTransposeA_CP_3763_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559/$exit
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612__entry__
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1501_to_assign_stmt_1559__exit__
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Update/cr
      -- 
    cr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1601_inst_req_1); -- 
    rr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1601_inst_req_0); -- 
    rr_4024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1585_inst_req_0); -- 
    cr_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1589_inst_req_1); -- 
    rr_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1589_inst_req_0); -- 
    cr_4029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1585_inst_req_1); -- 
    rr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1605_inst_req_0); -- 
    cr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(34), ack => type_cast_1605_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(23) & convTransposeA_CP_3763_elements(27) & convTransposeA_CP_3763_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Sample/ra
      -- 
    ra_4025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_0, ack => convTransposeA_CP_3763_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1585_Update/ca
      -- 
    ca_4030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_1, ack => convTransposeA_CP_3763_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_sample_completed_
      -- 
    ra_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_0, ack => convTransposeA_CP_3763_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1589_update_completed_
      -- 
    ca_4044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_1, ack => convTransposeA_CP_3763_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_sample_completed_
      -- 
    ra_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_0, ack => convTransposeA_CP_3763_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1601_update_completed_
      -- 
    ca_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_1, ack => convTransposeA_CP_3763_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Sample/ra
      -- 
    ra_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1605_inst_ack_0, ack => convTransposeA_CP_3763_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/type_cast_1605_Update/ca
      -- 
    ca_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1605_inst_ack_1, ack => convTransposeA_CP_3763_elements(42)); -- 
    -- CP-element group 43:  join  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (10) 
      -- CP-element group 43: 	 branch_block_stmt_1498/do_while_stmt_1636__entry__
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1498/merge_stmt_1614__exit__
      -- CP-element group 43: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612__exit__
      -- CP-element group 43: 	 branch_block_stmt_1498/assign_stmt_1566_to_assign_stmt_1612/$exit
      -- CP-element group 43: 	 branch_block_stmt_1498/merge_stmt_1614_PhiReqMerge
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/entry_whilex_xbody_PhiReq/$exit
      -- CP-element group 43: 	 branch_block_stmt_1498/merge_stmt_1614_PhiAck/$entry
      -- CP-element group 43: 	 branch_block_stmt_1498/merge_stmt_1614_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(36) & convTransposeA_CP_3763_elements(38) & convTransposeA_CP_3763_elements(40) & convTransposeA_CP_3763_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1498/do_while_stmt_1636/$entry
      -- CP-element group 44: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636__entry__
      -- 
    convTransposeA_CP_3763_elements(44) <= convTransposeA_CP_3763_elements(43);
    -- CP-element group 45:  merge  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	218 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636__exit__
      -- 
    -- Element group convTransposeA_CP_3763_elements(45) is bound as output of CP function.
    -- CP-element group 46:  merge  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_back
      -- 
    -- Element group convTransposeA_CP_3763_elements(46) is bound as output of CP function.
    -- CP-element group 47:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	52 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	217 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_taken/$entry
      -- CP-element group 47: 	 branch_block_stmt_1498/do_while_stmt_1636/condition_done
      -- CP-element group 47: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_exit/$entry
      -- 
    convTransposeA_CP_3763_elements(47) <= convTransposeA_CP_3763_elements(52);
    -- CP-element group 48:  branch  place  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	215 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_body_done
      -- 
    convTransposeA_CP_3763_elements(48) <= convTransposeA_CP_3763_elements(215);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	61 
    -- CP-element group 49: 	82 
    -- CP-element group 49: 	103 
    -- CP-element group 49: 	124 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/back_edge_to_loop_body
      -- 
    convTransposeA_CP_3763_elements(49) <= convTransposeA_CP_3763_elements(46);
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	44 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	63 
    -- CP-element group 50: 	84 
    -- CP-element group 50: 	105 
    -- CP-element group 50: 	126 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/first_time_through_loop_body
      -- 
    convTransposeA_CP_3763_elements(50) <= convTransposeA_CP_3763_elements(44);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	57 
    -- CP-element group 51: 	58 
    -- CP-element group 51: 	76 
    -- CP-element group 51: 	77 
    -- CP-element group 51: 	214 
    -- CP-element group 51: 	97 
    -- CP-element group 51: 	98 
    -- CP-element group 51: 	118 
    -- CP-element group 51: 	119 
    -- CP-element group 51: 	156 
    -- CP-element group 51: 	157 
    -- CP-element group 51: 	167 
    -- CP-element group 51: 	169 
    -- CP-element group 51: 	186 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/$entry
      -- CP-element group 51: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/loop_body_start
      -- 
    -- Element group convTransposeA_CP_3763_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	213 
    -- CP-element group 52: 	214 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	47 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/condition_evaluated
      -- 
    condition_evaluated_4087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(52), ack => do_while_stmt_1636_branch_req_0); -- 
    convTransposeA_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(56) & convTransposeA_CP_3763_elements(213) & convTransposeA_CP_3763_elements(214);
      gj_convTransposeA_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	57 
    -- CP-element group 53: 	76 
    -- CP-element group 53: 	97 
    -- CP-element group 53: 	118 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53: 	99 
    -- CP-element group 53: 	120 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/aggregated_phi_sample_req
      -- CP-element group 53: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_sample_start__ps
      -- 
    convTransposeA_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(57) & convTransposeA_CP_3763_elements(76) & convTransposeA_CP_3763_elements(97) & convTransposeA_CP_3763_elements(118) & convTransposeA_CP_3763_elements(56);
      gj_convTransposeA_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	59 
    -- CP-element group 54: 	79 
    -- CP-element group 54: 	100 
    -- CP-element group 54: 	121 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	207 
    -- CP-element group 54: 	215 
    -- CP-element group 54: 	195 
    -- CP-element group 54: 	199 
    -- CP-element group 54: 	203 
    -- CP-element group 54: 	183 
    -- CP-element group 54: 	187 
    -- CP-element group 54: 	191 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: 	76 
    -- CP-element group 54: 	97 
    -- CP-element group 54: 	118 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/aggregated_phi_sample_ack
      -- CP-element group 54: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_sample_completed_
      -- 
    convTransposeA_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(59) & convTransposeA_CP_3763_elements(79) & convTransposeA_CP_3763_elements(100) & convTransposeA_CP_3763_elements(121);
      gj_convTransposeA_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	77 
    -- CP-element group 55: 	98 
    -- CP-element group 55: 	119 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	80 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	122 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/aggregated_phi_update_req
      -- CP-element group 55: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_update_start__ps
      -- 
    convTransposeA_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(58) & convTransposeA_CP_3763_elements(77) & convTransposeA_CP_3763_elements(98) & convTransposeA_CP_3763_elements(119);
      gj_convTransposeA_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	81 
    -- CP-element group 56: 	102 
    -- CP-element group 56: 	123 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/aggregated_phi_update_ack
      -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(60) & convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(102) & convTransposeA_CP_3763_elements(123);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	53 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_sample_start_
      -- 
    convTransposeA_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(54);
      gj_convTransposeA_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	153 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	55 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_update_start_
      -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(60) & convTransposeA_CP_3763_elements(153);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: 	151 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	49 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_loopback_trigger
      -- 
    convTransposeA_CP_3763_elements(61) <= convTransposeA_CP_3763_elements(49);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_loopback_sample_req_ps
      -- 
    phi_stmt_1638_loopback_sample_req_4102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1638_loopback_sample_req_4102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(62), ack => phi_stmt_1638_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	50 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_entry_trigger
      -- 
    convTransposeA_CP_3763_elements(63) <= convTransposeA_CP_3763_elements(50);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_entry_sample_req_ps
      -- 
    phi_stmt_1638_entry_sample_req_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1638_entry_sample_req_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(64), ack => phi_stmt_1638_req_1); -- 
    -- Element group convTransposeA_CP_3763_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1638_phi_mux_ack_ps
      -- 
    phi_stmt_1638_phi_mux_ack_4108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1638_ack_0, ack => convTransposeA_CP_3763_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Sample/rr
      -- 
    rr_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(68), ack => type_cast_1641_inst_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(66) & convTransposeA_CP_3763_elements(70);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_update_start_
      -- CP-element group 69: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Update/cr
      -- 
    cr_4126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(69), ack => type_cast_1641_inst_req_1); -- 
    convTransposeA_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(67) & convTransposeA_CP_3763_elements(71);
      gj_convTransposeA_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Sample/ra
      -- 
    ra_4122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1641_inst_ack_0, ack => convTransposeA_CP_3763_elements(70)); -- 
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1641_Update/ca
      -- 
    ca_4127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1641_inst_ack_1, ack => convTransposeA_CP_3763_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_update_start_
      -- 
    -- Element group convTransposeA_CP_3763_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_update_completed__ps
      -- 
    convTransposeA_CP_3763_elements(74) <= convTransposeA_CP_3763_elements(75);
    -- CP-element group 75:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_indvar_at_entry_1642_update_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(73), ack => convTransposeA_CP_3763_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	51 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	54 
    -- CP-element group 76: 	193 
    -- CP-element group 76: 	185 
    -- CP-element group 76: 	189 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	53 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_sample_start_
      -- 
    convTransposeA_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(193) & convTransposeA_CP_3763_elements(185) & convTransposeA_CP_3763_elements(189);
      gj_convTransposeA_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	51 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: 	141 
    -- CP-element group 77: 	184 
    -- CP-element group 77: 	192 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	55 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_update_start_
      -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(141) & convTransposeA_CP_3763_elements(184) & convTransposeA_CP_3763_elements(192);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	53 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_sample_start__ps
      -- 
    convTransposeA_CP_3763_elements(78) <= convTransposeA_CP_3763_elements(53);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	54 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	55 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_update_start__ps
      -- 
    convTransposeA_CP_3763_elements(80) <= convTransposeA_CP_3763_elements(55);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	56 
    -- CP-element group 81: 	139 
    -- CP-element group 81: 	182 
    -- CP-element group 81: 	190 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	49 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_loopback_trigger
      -- 
    convTransposeA_CP_3763_elements(82) <= convTransposeA_CP_3763_elements(49);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_loopback_sample_req_ps
      -- 
    phi_stmt_1643_loopback_sample_req_4146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1643_loopback_sample_req_4146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(83), ack => phi_stmt_1643_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	50 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_entry_trigger
      -- 
    convTransposeA_CP_3763_elements(84) <= convTransposeA_CP_3763_elements(50);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_entry_sample_req_ps
      -- 
    phi_stmt_1643_entry_sample_req_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1643_entry_sample_req_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(85), ack => phi_stmt_1643_req_1); -- 
    -- Element group convTransposeA_CP_3763_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_phi_mux_ack
      -- CP-element group 86: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1643_phi_mux_ack_ps
      -- 
    phi_stmt_1643_phi_mux_ack_4152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1643_ack_0, ack => convTransposeA_CP_3763_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Sample/rr
      -- 
    rr_4165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(89), ack => type_cast_1646_inst_req_0); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(87) & convTransposeA_CP_3763_elements(91);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_update_start_
      -- CP-element group 90: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Update/cr
      -- 
    cr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(90), ack => type_cast_1646_inst_req_1); -- 
    convTransposeA_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(88) & convTransposeA_CP_3763_elements(92);
      gj_convTransposeA_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Sample/ra
      -- 
    ra_4166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_0, ack => convTransposeA_CP_3763_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1646_Update/ca
      -- 
    ca_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_1, ack => convTransposeA_CP_3763_elements(92)); -- 
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_sample_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_update_start_
      -- 
    -- Element group convTransposeA_CP_3763_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_update_completed__ps
      -- 
    convTransposeA_CP_3763_elements(95) <= convTransposeA_CP_3763_elements(96);
    -- CP-element group 96:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim2x_x1_at_entry_1647_update_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(94), ack => convTransposeA_CP_3763_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	51 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	54 
    -- CP-element group 97: 	197 
    -- CP-element group 97: 	201 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	53 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_sample_start_
      -- 
    convTransposeA_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(197) & convTransposeA_CP_3763_elements(201);
      gj_convTransposeA_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	51 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: 	145 
    -- CP-element group 98: 	200 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	55 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_update_start_
      -- 
    convTransposeA_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(102) & convTransposeA_CP_3763_elements(145) & convTransposeA_CP_3763_elements(200);
      gj_convTransposeA_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	53 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_sample_start__ps
      -- 
    convTransposeA_CP_3763_elements(99) <= convTransposeA_CP_3763_elements(53);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	54 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_update_start__ps
      -- 
    convTransposeA_CP_3763_elements(101) <= convTransposeA_CP_3763_elements(55);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	56 
    -- CP-element group 102: 	143 
    -- CP-element group 102: 	198 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	49 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_loopback_trigger
      -- 
    convTransposeA_CP_3763_elements(103) <= convTransposeA_CP_3763_elements(49);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_loopback_sample_req_ps
      -- 
    phi_stmt_1648_loopback_sample_req_4190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1648_loopback_sample_req_4190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(104), ack => phi_stmt_1648_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	50 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_entry_trigger
      -- 
    convTransposeA_CP_3763_elements(105) <= convTransposeA_CP_3763_elements(50);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_entry_sample_req_ps
      -- 
    phi_stmt_1648_entry_sample_req_4193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1648_entry_sample_req_4193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(106), ack => phi_stmt_1648_req_1); -- 
    -- Element group convTransposeA_CP_3763_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1648_phi_mux_ack_ps
      -- 
    phi_stmt_1648_phi_mux_ack_4196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1648_ack_0, ack => convTransposeA_CP_3763_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Sample/rr
      -- 
    rr_4209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(110), ack => type_cast_1651_inst_req_0); -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(108) & convTransposeA_CP_3763_elements(112);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Update/cr
      -- 
    cr_4214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(111), ack => type_cast_1651_inst_req_1); -- 
    convTransposeA_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(109) & convTransposeA_CP_3763_elements(113);
      gj_convTransposeA_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Sample/ra
      -- 
    ra_4210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_0, ack => convTransposeA_CP_3763_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1651_Update/ca
      -- 
    ca_4215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_1, ack => convTransposeA_CP_3763_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_update_start_
      -- 
    -- Element group convTransposeA_CP_3763_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_update_completed__ps
      -- 
    convTransposeA_CP_3763_elements(116) <= convTransposeA_CP_3763_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim1x_x1_at_entry_1652_update_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(115), ack => convTransposeA_CP_3763_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	51 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	54 
    -- CP-element group 118: 	205 
    -- CP-element group 118: 	209 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	53 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_sample_start_
      -- 
    convTransposeA_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(205) & convTransposeA_CP_3763_elements(209);
      gj_convTransposeA_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	51 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	208 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	149 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	55 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_update_start_
      -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(208) & convTransposeA_CP_3763_elements(123) & convTransposeA_CP_3763_elements(149);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	53 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_sample_start__ps
      -- 
    convTransposeA_CP_3763_elements(120) <= convTransposeA_CP_3763_elements(53);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	54 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_sample_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	55 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_update_start__ps
      -- 
    convTransposeA_CP_3763_elements(122) <= convTransposeA_CP_3763_elements(55);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	56 
    -- CP-element group 123: 	206 
    -- CP-element group 123: 	147 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	119 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_update_completed__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	49 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_loopback_trigger
      -- 
    convTransposeA_CP_3763_elements(124) <= convTransposeA_CP_3763_elements(49);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_loopback_sample_req
      -- CP-element group 125: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_loopback_sample_req_ps
      -- 
    phi_stmt_1653_loopback_sample_req_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1653_loopback_sample_req_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(125), ack => phi_stmt_1653_req_0); -- 
    -- Element group convTransposeA_CP_3763_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	50 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_entry_trigger
      -- 
    convTransposeA_CP_3763_elements(126) <= convTransposeA_CP_3763_elements(50);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_entry_sample_req_ps
      -- 
    phi_stmt_1653_entry_sample_req_4237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1653_entry_sample_req_4237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(127), ack => phi_stmt_1653_req_1); -- 
    -- Element group convTransposeA_CP_3763_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_phi_mux_ack_ps
      -- CP-element group 128: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/phi_stmt_1653_phi_mux_ack
      -- 
    phi_stmt_1653_phi_mux_ack_4240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1653_ack_0, ack => convTransposeA_CP_3763_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_sample_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_update_start__ps
      -- 
    -- Element group convTransposeA_CP_3763_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Sample/rr
      -- 
    rr_4253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(131), ack => type_cast_1656_inst_req_0); -- 
    convTransposeA_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(129) & convTransposeA_CP_3763_elements(133);
      gj_convTransposeA_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_update_start_
      -- CP-element group 132: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Update/cr
      -- 
    cr_4258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(132), ack => type_cast_1656_inst_req_1); -- 
    convTransposeA_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(130) & convTransposeA_CP_3763_elements(134);
      gj_convTransposeA_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Sample/ra
      -- 
    ra_4254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1656_inst_ack_0, ack => convTransposeA_CP_3763_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1656_Update/ca
      -- 
    ca_4259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1656_inst_ack_1, ack => convTransposeA_CP_3763_elements(134)); -- 
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_sample_start__ps
      -- CP-element group 135: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_sample_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_update_start__ps
      -- CP-element group 136: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_update_start_
      -- 
    -- Element group convTransposeA_CP_3763_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_update_completed__ps
      -- 
    convTransposeA_CP_3763_elements(137) <= convTransposeA_CP_3763_elements(138);
    -- CP-element group 138:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	137 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/R_input_dim0x_x1_at_entry_1657_update_completed_
      -- 
    -- Element group convTransposeA_CP_3763_elements(138) is a control-delay.
    cp_element_138_delay: control_delay_element  generic map(name => " 138_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(136), ack => convTransposeA_CP_3763_elements(138), clk => clk, reset =>reset);
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	81 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Sample/rr
      -- 
    rr_4276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(139), ack => type_cast_1686_inst_req_0); -- 
    convTransposeA_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(141);
      gj_convTransposeA_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: 	170 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_update_start_
      -- CP-element group 140: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Update/cr
      -- 
    cr_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(140), ack => type_cast_1686_inst_req_1); -- 
    convTransposeA_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(142) & convTransposeA_CP_3763_elements(170);
      gj_convTransposeA_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	77 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Sample/ra
      -- 
    ra_4277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_0, ack => convTransposeA_CP_3763_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	168 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1686_Update/ca
      -- 
    ca_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_1, ack => convTransposeA_CP_3763_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	102 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Sample/rr
      -- 
    rr_4290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(143), ack => type_cast_1690_inst_req_0); -- 
    convTransposeA_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(102) & convTransposeA_CP_3763_elements(145);
      gj_convTransposeA_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: 	170 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Update/cr
      -- 
    cr_4295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(144), ack => type_cast_1690_inst_req_1); -- 
    convTransposeA_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(146) & convTransposeA_CP_3763_elements(170);
      gj_convTransposeA_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	98 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Sample/ra
      -- 
    ra_4291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1690_inst_ack_0, ack => convTransposeA_CP_3763_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	168 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1690_Update/ca
      -- 
    ca_4296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1690_inst_ack_1, ack => convTransposeA_CP_3763_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	123 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Sample/rr
      -- 
    rr_4304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(147), ack => type_cast_1694_inst_req_0); -- 
    convTransposeA_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(123) & convTransposeA_CP_3763_elements(149);
      gj_convTransposeA_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: 	170 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_update_start_
      -- CP-element group 148: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Update/cr
      -- 
    cr_4309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(148), ack => type_cast_1694_inst_req_1); -- 
    convTransposeA_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(150) & convTransposeA_CP_3763_elements(170);
      gj_convTransposeA_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	119 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Sample/ra
      -- 
    ra_4305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_0, ack => convTransposeA_CP_3763_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	168 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1694_Update/ca
      -- 
    ca_4310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1694_inst_ack_1, ack => convTransposeA_CP_3763_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	60 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Sample/rr
      -- 
    rr_4318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(151), ack => type_cast_1718_inst_req_0); -- 
    convTransposeA_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(60) & convTransposeA_CP_3763_elements(153);
      gj_convTransposeA_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: 	158 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_update_start_
      -- CP-element group 152: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Update/cr
      -- 
    cr_4323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(152), ack => type_cast_1718_inst_req_1); -- 
    convTransposeA_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(154) & convTransposeA_CP_3763_elements(158);
      gj_convTransposeA_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	58 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Sample/ra
      -- 
    ra_4319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_0, ack => convTransposeA_CP_3763_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	158 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (16) 
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1718_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_resized_1
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_scaled_1
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_computed_1
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_resize_1/$entry
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_resize_1/$exit
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_resize_1/index_resize_req
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_resize_1/index_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_scale_1/$entry
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_scale_1/$exit
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_scale_1/scale_rename_req
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_index_scale_1/scale_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Sample/req
      -- 
    ca_4324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_1, ack => convTransposeA_CP_3763_elements(154)); -- 
    req_4349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(154), ack => array_obj_ref_1724_index_offset_req_0); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	160 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	160 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_request/$entry
      -- CP-element group 155: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_request/req
      -- 
    req_4364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(155), ack => addr_of_1725_final_reg_req_0); -- 
    convTransposeA_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(159) & convTransposeA_CP_3763_elements(160);
      gj_convTransposeA_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	51 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	164 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_update_start_
      -- CP-element group 156: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_complete/req
      -- 
    req_4369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(156), ack => addr_of_1725_final_reg_req_1); -- 
    convTransposeA_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(161) & convTransposeA_CP_3763_elements(164);
      gj_convTransposeA_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	51 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_update_start
      -- CP-element group 157: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Update/req
      -- 
    req_4354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(157), ack => array_obj_ref_1724_index_offset_req_1); -- 
    convTransposeA_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(159) & convTransposeA_CP_3763_elements(160);
      gj_convTransposeA_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	215 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	152 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_sample_complete
      -- CP-element group 158: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Sample/ack
      -- 
    ack_4350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1724_index_offset_ack_0, ack => convTransposeA_CP_3763_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (8) 
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_root_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_offset_calculated
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_final_index_sum_regn_Update/ack
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_base_plus_offset/$entry
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_base_plus_offset/$exit
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_base_plus_offset/sum_rename_req
      -- CP-element group 159: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1724_base_plus_offset/sum_rename_ack
      -- 
    ack_4355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1724_index_offset_ack_1, ack => convTransposeA_CP_3763_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_request/$exit
      -- CP-element group 160: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_request/ack
      -- 
    ack_4365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1725_final_reg_ack_0, ack => convTransposeA_CP_3763_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (19) 
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_complete/$exit
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1725_complete/ack
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_word_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_root_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_address_resized
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_addr_resize/$entry
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_addr_resize/$exit
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_addr_resize/base_resize_req
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_addr_resize/base_resize_ack
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_plus_offset/$entry
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_plus_offset/$exit
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_plus_offset/sum_rename_req
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_base_plus_offset/sum_rename_ack
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_word_addrgen/$entry
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_word_addrgen/$exit
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_word_addrgen/root_register_req
      -- CP-element group 161: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_word_addrgen/root_register_ack
      -- 
    ack_4370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1725_final_reg_ack_1, ack => convTransposeA_CP_3763_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/word_access_start/word_0/rr
      -- CP-element group 162: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/word_access_start/word_0/$entry
      -- 
    rr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(162), ack => ptr_deref_1729_load_0_req_0); -- 
    convTransposeA_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(161) & convTransposeA_CP_3763_elements(164);
      gj_convTransposeA_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: 	180 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_update_start_
      -- 
    cr_4414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(163), ack => ptr_deref_1729_load_0_req_1); -- 
    convTransposeA_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(165) & convTransposeA_CP_3763_elements(180);
      gj_convTransposeA_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/word_access_start/word_0/ra
      -- CP-element group 164: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/word_access_start/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Sample/word_access_start/$exit
      -- 
    ra_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1729_load_0_ack_0, ack => convTransposeA_CP_3763_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	178 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (9) 
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/word_access_complete/word_0/ca
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/word_access_complete/word_0/$exit
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/ptr_deref_1729_Merge/$entry
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/word_access_complete/$exit
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/ptr_deref_1729_Merge/merge_ack
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/ptr_deref_1729_Merge/merge_req
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_Update/ptr_deref_1729_Merge/$exit
      -- CP-element group 165: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1729_update_completed_
      -- 
    ca_4415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1729_load_0_ack_1, ack => convTransposeA_CP_3763_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	171 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	172 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	172 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_request/$entry
      -- CP-element group 166: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_request/req
      -- 
    req_4460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(166), ack => addr_of_1748_final_reg_req_0); -- 
    convTransposeA_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(171) & convTransposeA_CP_3763_elements(172);
      gj_convTransposeA_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	51 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	173 
    -- CP-element group 167: 	176 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	173 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_complete/req
      -- CP-element group 167: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_update_start_
      -- CP-element group 167: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_complete/$entry
      -- 
    req_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(167), ack => addr_of_1748_final_reg_req_1); -- 
    convTransposeA_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(173) & convTransposeA_CP_3763_elements(176);
      gj_convTransposeA_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	142 
    -- CP-element group 168: 	146 
    -- CP-element group 168: 	150 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (13) 
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_resized_1
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Sample/req
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_scale_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_scale_1/scale_rename_req
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_scale_1/scale_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_scale_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_resize_1/index_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_resize_1/index_resize_req
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_resize_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_resize_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_computed_1
      -- CP-element group 168: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_index_scaled_1
      -- 
    req_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(168), ack => array_obj_ref_1747_index_offset_req_0); -- 
    convTransposeA_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(142) & convTransposeA_CP_3763_elements(146) & convTransposeA_CP_3763_elements(150);
      gj_convTransposeA_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	51 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_update_start
      -- CP-element group 169: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Update/req
      -- 
    req_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(169), ack => array_obj_ref_1747_index_offset_req_1); -- 
    convTransposeA_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(171) & convTransposeA_CP_3763_elements(172);
      gj_convTransposeA_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	215 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	140 
    -- CP-element group 170: 	144 
    -- CP-element group 170: 	148 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Sample/ack
      -- CP-element group 170: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_sample_complete
      -- 
    ack_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1747_index_offset_ack_0, ack => convTransposeA_CP_3763_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	166 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (8) 
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/array_obj_ref_1747_base_plus_offset/sum_rename_ack
      -- 
    ack_4451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1747_index_offset_ack_1, ack => convTransposeA_CP_3763_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_request/ack
      -- CP-element group 172: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_request/$exit
      -- 
    ack_4461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1748_final_reg_ack_0, ack => convTransposeA_CP_3763_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	167 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	167 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_complete/ack
      -- CP-element group 173: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/addr_of_1748_complete/$exit
      -- 
    ack_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1748_final_reg_ack_1, ack => convTransposeA_CP_3763_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Sample/req
      -- CP-element group 174: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Sample/$entry
      -- 
    req_4474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(174), ack => W_arrayidx81_1750_delayed_6_0_1750_inst_req_0); -- 
    convTransposeA_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(173) & convTransposeA_CP_3763_elements(176);
      gj_convTransposeA_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: 	180 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Update/req
      -- CP-element group 175: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Update/$entry
      -- 
    req_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(175), ack => W_arrayidx81_1750_delayed_6_0_1750_inst_req_1); -- 
    convTransposeA_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(177) & convTransposeA_CP_3763_elements(180);
      gj_convTransposeA_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	167 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Sample/ack
      -- CP-element group 176: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Sample/$exit
      -- 
    ack_4475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx81_1750_delayed_6_0_1750_inst_ack_0, ack => convTransposeA_CP_3763_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (19) 
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_word_addrgen/root_register_ack
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_word_addrgen/root_register_req
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_word_addrgen/$exit
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_word_addrgen/$entry
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_plus_offset/sum_rename_ack
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_plus_offset/sum_rename_req
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_plus_offset/$exit
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_plus_offset/$entry
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_addr_resize/base_resize_ack
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_addr_resize/base_resize_req
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_addr_resize/$exit
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_addr_resize/$entry
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_address_resized
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_root_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_word_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_base_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Update/ack
      -- CP-element group 177: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1752_Update/$exit
      -- 
    ack_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx81_1750_delayed_6_0_1750_inst_ack_1, ack => convTransposeA_CP_3763_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	165 
    -- CP-element group 178: 	177 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/word_access_start/word_0/$entry
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/word_access_start/$entry
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/ptr_deref_1754_Split/split_ack
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/word_access_start/word_0/rr
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/ptr_deref_1754_Split/split_req
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/ptr_deref_1754_Split/$exit
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/ptr_deref_1754_Split/$entry
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_sample_start_
      -- 
    rr_4518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(178), ack => ptr_deref_1754_store_0_req_0); -- 
    convTransposeA_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(165) & convTransposeA_CP_3763_elements(177) & convTransposeA_CP_3763_elements(180);
      gj_convTransposeA_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (5) 
      -- CP-element group 179: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/word_access_complete/$entry
      -- CP-element group 179: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/word_access_complete/word_0/cr
      -- CP-element group 179: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/word_access_complete/word_0/$entry
      -- CP-element group 179: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_update_start_
      -- 
    cr_4529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(179), ack => ptr_deref_1754_store_0_req_1); -- 
    convTransposeA_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeA_CP_3763_elements(181);
      gj_convTransposeA_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	163 
    -- CP-element group 180: 	175 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/word_access_start/$exit
      -- CP-element group 180: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/word_access_start/word_0/$exit
      -- CP-element group 180: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/word_access_start/word_0/ra
      -- CP-element group 180: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_sample_completed_
      -- 
    ra_4519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1754_store_0_ack_0, ack => convTransposeA_CP_3763_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	215 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/word_access_complete/word_0/ca
      -- CP-element group 181: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/word_access_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_Update/word_access_complete/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/ptr_deref_1754_update_completed_
      -- 
    ca_4530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1754_store_0_ack_1, ack => convTransposeA_CP_3763_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	81 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Sample/rr
      -- 
    rr_4538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(182), ack => type_cast_1759_inst_req_0); -- 
    convTransposeA_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(184);
      gj_convTransposeA_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	54 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	196 
    -- CP-element group 183: 	185 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Update/cr
      -- 
    cr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(183), ack => type_cast_1759_inst_req_1); -- 
    convTransposeA_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(196) & convTransposeA_CP_3763_elements(185);
      gj_convTransposeA_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	77 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Sample/ra
      -- CP-element group 184: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_sample_completed_
      -- 
    ra_4539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_0, ack => convTransposeA_CP_3763_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	194 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	76 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1759_update_completed_
      -- 
    ca_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_1, ack => convTransposeA_CP_3763_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	51 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Sample/$entry
      -- 
    rr_4552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(186), ack => type_cast_1763_inst_req_0); -- 
    convTransposeA_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(51) & convTransposeA_CP_3763_elements(188);
      gj_convTransposeA_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	54 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	196 
    -- CP-element group 187: 	189 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Update/$entry
      -- 
    cr_4557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(187), ack => type_cast_1763_inst_req_1); -- 
    convTransposeA_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(196) & convTransposeA_CP_3763_elements(189);
      gj_convTransposeA_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Sample/ra
      -- 
    ra_4553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1763_inst_ack_0, ack => convTransposeA_CP_3763_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	194 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	76 
    -- CP-element group 189: 	187 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1763_update_completed_
      -- 
    ca_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1763_inst_ack_1, ack => convTransposeA_CP_3763_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	81 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Sample/req
      -- CP-element group 190: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Sample/$entry
      -- 
    req_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(190), ack => W_add96_1773_delayed_1_0_1777_inst_req_0); -- 
    convTransposeA_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(81) & convTransposeA_CP_3763_elements(192);
      gj_convTransposeA_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	54 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Update/req
      -- CP-element group 191: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_update_start_
      -- 
    req_4571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(191), ack => W_add96_1773_delayed_1_0_1777_inst_req_1); -- 
    convTransposeA_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(193);
      gj_convTransposeA_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	77 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Sample/ack
      -- CP-element group 192: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_sample_completed_
      -- 
    ack_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add96_1773_delayed_1_0_1777_inst_ack_0, ack => convTransposeA_CP_3763_elements(192)); -- 
    -- CP-element group 193:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	215 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	76 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Update/ack
      -- CP-element group 193: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1779_update_completed_
      -- 
    ack_4572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add96_1773_delayed_1_0_1777_inst_ack_1, ack => convTransposeA_CP_3763_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	185 
    -- CP-element group 194: 	189 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_sample_start_
      -- 
    rr_4580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(194), ack => type_cast_1789_inst_req_0); -- 
    convTransposeA_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(185) & convTransposeA_CP_3763_elements(189) & convTransposeA_CP_3763_elements(196);
      gj_convTransposeA_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	54 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	204 
    -- CP-element group 195: 	197 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Update/cr
      -- 
    cr_4585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(195), ack => type_cast_1789_inst_req_1); -- 
    convTransposeA_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(204) & convTransposeA_CP_3763_elements(197);
      gj_convTransposeA_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: 	183 
    -- CP-element group 196: 	187 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Sample/ra
      -- CP-element group 196: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_sample_completed_
      -- 
    ra_4581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1789_inst_ack_0, ack => convTransposeA_CP_3763_elements(196)); -- 
    -- CP-element group 197:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	202 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	97 
    -- CP-element group 197: 	195 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1789_Update/ca
      -- 
    ca_4586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1789_inst_ack_1, ack => convTransposeA_CP_3763_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	102 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Sample/req
      -- 
    req_4594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(198), ack => W_input_dim1x_x1_1790_delayed_2_0_1797_inst_req_0); -- 
    convTransposeA_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(102) & convTransposeA_CP_3763_elements(200);
      gj_convTransposeA_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	54 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	204 
    -- CP-element group 199: 	201 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Update/req
      -- CP-element group 199: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_update_start_
      -- 
    req_4599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(199), ack => W_input_dim1x_x1_1790_delayed_2_0_1797_inst_req_1); -- 
    convTransposeA_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(204) & convTransposeA_CP_3763_elements(201);
      gj_convTransposeA_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	98 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Sample/ack
      -- CP-element group 200: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_sample_completed_
      -- 
    ack_4595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_1790_delayed_2_0_1797_inst_ack_0, ack => convTransposeA_CP_3763_elements(200)); -- 
    -- CP-element group 201:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	97 
    -- CP-element group 201: 	199 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1799_Update/ack
      -- 
    ack_4600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_1790_delayed_2_0_1797_inst_ack_1, ack => convTransposeA_CP_3763_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	197 
    -- CP-element group 202: 	201 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Sample/rr
      -- 
    rr_4608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(202), ack => type_cast_1812_inst_req_0); -- 
    convTransposeA_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(197) & convTransposeA_CP_3763_elements(201) & convTransposeA_CP_3763_elements(204);
      gj_convTransposeA_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	54 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: 	212 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_update_start_
      -- CP-element group 203: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Update/cr
      -- CP-element group 203: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Update/$entry
      -- 
    cr_4613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(203), ack => type_cast_1812_inst_req_1); -- 
    convTransposeA_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(205) & convTransposeA_CP_3763_elements(212);
      gj_convTransposeA_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	195 
    -- CP-element group 204: 	199 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Sample/$exit
      -- 
    ra_4609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1812_inst_ack_0, ack => convTransposeA_CP_3763_elements(204)); -- 
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	210 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	118 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1812_Update/$exit
      -- 
    ca_4614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1812_inst_ack_1, ack => convTransposeA_CP_3763_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	123 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Sample/req
      -- 
    req_4622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(206), ack => W_input_dim0x_x1_1804_delayed_3_0_1814_inst_req_0); -- 
    convTransposeA_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(123) & convTransposeA_CP_3763_elements(208);
      gj_convTransposeA_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	54 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: 	212 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_update_start_
      -- CP-element group 207: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Update/req
      -- CP-element group 207: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Update/$entry
      -- 
    req_4627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(207), ack => W_input_dim0x_x1_1804_delayed_3_0_1814_inst_req_1); -- 
    convTransposeA_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(209) & convTransposeA_CP_3763_elements(212);
      gj_convTransposeA_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: 	119 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Sample/ack
      -- 
    ack_4623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_1804_delayed_3_0_1814_inst_ack_0, ack => convTransposeA_CP_3763_elements(208)); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: 	118 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Update/ack
      -- CP-element group 209: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/assign_stmt_1816_Update/$exit
      -- 
    ack_4628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_1804_delayed_3_0_1814_inst_ack_1, ack => convTransposeA_CP_3763_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	205 
    -- CP-element group 210: 	209 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Sample/rr
      -- 
    rr_4636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(210), ack => type_cast_1831_inst_req_0); -- 
    convTransposeA_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(205) & convTransposeA_CP_3763_elements(209) & convTransposeA_CP_3763_elements(212);
      gj_convTransposeA_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_update_start_
      -- CP-element group 211: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Update/$entry
      -- 
    cr_4641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(211), ack => type_cast_1831_inst_req_1); -- 
    convTransposeA_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeA_CP_3763_elements(213);
      gj_convTransposeA_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	207 
    -- CP-element group 212: 	210 
    -- CP-element group 212: 	203 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Sample/ra
      -- CP-element group 212: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Sample/$exit
      -- 
    ra_4637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_0, ack => convTransposeA_CP_3763_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	52 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/type_cast_1831_Update/$exit
      -- 
    ca_4642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_1, ack => convTransposeA_CP_3763_elements(213)); -- 
    -- CP-element group 214:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	51 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	52 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convTransposeA_CP_3763_elements(214) is a control-delay.
    cp_element_214_delay: control_delay_element  generic map(name => " 214_delay", delay_value => 1)  port map(req => convTransposeA_CP_3763_elements(51), ack => convTransposeA_CP_3763_elements(214), clk => clk, reset =>reset);
    -- CP-element group 215:  join  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	54 
    -- CP-element group 215: 	158 
    -- CP-element group 215: 	170 
    -- CP-element group 215: 	193 
    -- CP-element group 215: 	181 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	48 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_1498/do_while_stmt_1636/do_while_stmt_1636_loop_body/$exit
      -- 
    convTransposeA_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeA_CP_3763_elements(54) & convTransposeA_CP_3763_elements(158) & convTransposeA_CP_3763_elements(170) & convTransposeA_CP_3763_elements(193) & convTransposeA_CP_3763_elements(181);
      gj_convTransposeA_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3763_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_exit/ack
      -- CP-element group 216: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_exit/$exit
      -- 
    ack_4647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1636_branch_ack_0, ack => convTransposeA_CP_3763_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	47 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_taken/ack
      -- CP-element group 217: 	 branch_block_stmt_1498/do_while_stmt_1636/loop_taken/$exit
      -- 
    ack_4651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1636_branch_ack_1, ack => convTransposeA_CP_3763_elements(217)); -- 
    -- CP-element group 218:  transition  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	1 
    -- CP-element group 218:  members (1) 
      -- CP-element group 218: 	 branch_block_stmt_1498/do_while_stmt_1636/$exit
      -- 
    convTransposeA_CP_3763_elements(218) <= convTransposeA_CP_3763_elements(45);
    -- CP-element group 219:  merge  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	1 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (15) 
      -- CP-element group 219: 	 branch_block_stmt_1498/merge_stmt_1854__exit__
      -- CP-element group 219: 	 branch_block_stmt_1498/assign_stmt_1859__entry__
      -- CP-element group 219: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_1498/assign_stmt_1859/$entry
      -- CP-element group 219: 	 branch_block_stmt_1498/if_stmt_1850_if_link/if_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_1498/if_stmt_1850_if_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_1498/whilex_xbody_whilex_xend
      -- CP-element group 219: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_1498/merge_stmt_1854_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Sample/req
      -- CP-element group 219: 	 branch_block_stmt_1498/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_1498/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_1498/merge_stmt_1854_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_1498/merge_stmt_1854_PhiAck/$exit
      -- CP-element group 219: 	 branch_block_stmt_1498/merge_stmt_1854_PhiAck/dummy
      -- 
    if_choice_transition_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1850_branch_ack_1, ack => convTransposeA_CP_3763_elements(219)); -- 
    req_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(219), ack => WPIPE_Block0_done_1856_inst_req_0); -- 
    -- CP-element group 220:  merge  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	1 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_1498/if_stmt_1850__exit__
      -- CP-element group 220: 	 branch_block_stmt_1498/merge_stmt_1854__entry__
      -- CP-element group 220: 	 branch_block_stmt_1498/if_stmt_1850_else_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_1498/if_stmt_1850_else_link/else_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_1498/merge_stmt_1854_dead_link/$entry
      -- 
    else_choice_transition_4669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1850_branch_ack_0, ack => convTransposeA_CP_3763_elements(220)); -- 
    -- CP-element group 221:  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_update_start_
      -- CP-element group 221: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Sample/ack
      -- CP-element group 221: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Update/req
      -- 
    ack_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1856_inst_ack_0, ack => convTransposeA_CP_3763_elements(221)); -- 
    req_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3763_elements(221), ack => WPIPE_Block0_done_1856_inst_req_1); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (16) 
      -- CP-element group 222: 	 branch_block_stmt_1498/assign_stmt_1859__exit__
      -- CP-element group 222: 	 $exit
      -- CP-element group 222: 	 branch_block_stmt_1498/$exit
      -- CP-element group 222: 	 branch_block_stmt_1498/branch_block_stmt_1498__exit__
      -- CP-element group 222: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_1498/assign_stmt_1859/$exit
      -- CP-element group 222: 	 branch_block_stmt_1498/return__
      -- CP-element group 222: 	 branch_block_stmt_1498/merge_stmt_1861__exit__
      -- CP-element group 222: 	 branch_block_stmt_1498/merge_stmt_1861_PhiReqMerge
      -- CP-element group 222: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_1498/assign_stmt_1859/WPIPE_Block0_done_1856_Update/ack
      -- CP-element group 222: 	 branch_block_stmt_1498/return___PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_1498/return___PhiReq/$exit
      -- CP-element group 222: 	 branch_block_stmt_1498/merge_stmt_1861_PhiAck/$entry
      -- CP-element group 222: 	 branch_block_stmt_1498/merge_stmt_1861_PhiAck/$exit
      -- CP-element group 222: 	 branch_block_stmt_1498/merge_stmt_1861_PhiAck/dummy
      -- 
    ack_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1856_inst_ack_1, ack => convTransposeA_CP_3763_elements(222)); -- 
    convTransposeA_do_while_stmt_1636_terminator_4652: loop_terminator -- 
      generic map (name => " convTransposeA_do_while_stmt_1636_terminator_4652", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convTransposeA_CP_3763_elements(48),loop_continue => convTransposeA_CP_3763_elements(217),loop_terminate => convTransposeA_CP_3763_elements(216),loop_back => convTransposeA_CP_3763_elements(46),loop_exit => convTransposeA_CP_3763_elements(45),clk => clk, reset => reset); -- 
    phi_stmt_1638_phi_seq_4136_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3763_elements(61);
      convTransposeA_CP_3763_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3763_elements(70);
      convTransposeA_CP_3763_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3763_elements(71);
      convTransposeA_CP_3763_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3763_elements(63);
      convTransposeA_CP_3763_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3763_elements(72);
      convTransposeA_CP_3763_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3763_elements(74);
      convTransposeA_CP_3763_elements(64) <= phi_mux_reqs(1);
      phi_stmt_1638_phi_seq_4136 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1638_phi_seq_4136") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3763_elements(53), 
          phi_sample_ack => convTransposeA_CP_3763_elements(59), 
          phi_update_req => convTransposeA_CP_3763_elements(55), 
          phi_update_ack => convTransposeA_CP_3763_elements(60), 
          phi_mux_ack => convTransposeA_CP_3763_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1643_phi_seq_4180_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3763_elements(82);
      convTransposeA_CP_3763_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3763_elements(91);
      convTransposeA_CP_3763_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3763_elements(92);
      convTransposeA_CP_3763_elements(83) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3763_elements(84);
      convTransposeA_CP_3763_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3763_elements(93);
      convTransposeA_CP_3763_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3763_elements(95);
      convTransposeA_CP_3763_elements(85) <= phi_mux_reqs(1);
      phi_stmt_1643_phi_seq_4180 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1643_phi_seq_4180") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3763_elements(78), 
          phi_sample_ack => convTransposeA_CP_3763_elements(79), 
          phi_update_req => convTransposeA_CP_3763_elements(80), 
          phi_update_ack => convTransposeA_CP_3763_elements(81), 
          phi_mux_ack => convTransposeA_CP_3763_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1648_phi_seq_4224_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3763_elements(103);
      convTransposeA_CP_3763_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3763_elements(112);
      convTransposeA_CP_3763_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3763_elements(113);
      convTransposeA_CP_3763_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3763_elements(105);
      convTransposeA_CP_3763_elements(114)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3763_elements(114);
      convTransposeA_CP_3763_elements(115)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3763_elements(116);
      convTransposeA_CP_3763_elements(106) <= phi_mux_reqs(1);
      phi_stmt_1648_phi_seq_4224 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1648_phi_seq_4224") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3763_elements(99), 
          phi_sample_ack => convTransposeA_CP_3763_elements(100), 
          phi_update_req => convTransposeA_CP_3763_elements(101), 
          phi_update_ack => convTransposeA_CP_3763_elements(102), 
          phi_mux_ack => convTransposeA_CP_3763_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1653_phi_seq_4268_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeA_CP_3763_elements(124);
      convTransposeA_CP_3763_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeA_CP_3763_elements(133);
      convTransposeA_CP_3763_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeA_CP_3763_elements(134);
      convTransposeA_CP_3763_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeA_CP_3763_elements(126);
      convTransposeA_CP_3763_elements(135)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeA_CP_3763_elements(135);
      convTransposeA_CP_3763_elements(136)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeA_CP_3763_elements(137);
      convTransposeA_CP_3763_elements(127) <= phi_mux_reqs(1);
      phi_stmt_1653_phi_seq_4268 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1653_phi_seq_4268") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeA_CP_3763_elements(120), 
          phi_sample_ack => convTransposeA_CP_3763_elements(121), 
          phi_update_req => convTransposeA_CP_3763_elements(122), 
          phi_update_ack => convTransposeA_CP_3763_elements(123), 
          phi_mux_ack => convTransposeA_CP_3763_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4088_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convTransposeA_CP_3763_elements(49);
        preds(1)  <= convTransposeA_CP_3763_elements(50);
        entry_tmerge_4088 : transition_merge -- 
          generic map(name => " entry_tmerge_4088")
          port map (preds => preds, symbol_out => convTransposeA_CP_3763_elements(51));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_1849_wire : std_logic_vector(0 downto 0);
    signal R_idxprom80_1746_resized : std_logic_vector(13 downto 0);
    signal R_idxprom80_1746_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1723_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1723_scaled : std_logic_vector(13 downto 0);
    signal add41_1566 : std_logic_vector(15 downto 0);
    signal add54_1577 : std_logic_vector(15 downto 0);
    signal add73_1705 : std_logic_vector(63 downto 0);
    signal add75_1715 : std_logic_vector(63 downto 0);
    signal add96_1773_delayed_1_0_1779 : std_logic_vector(15 downto 0);
    signal add96_1776 : std_logic_vector(15 downto 0);
    signal add_1550 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1663 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1724_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1724_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1724_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1724_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1724_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1724_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1747_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1747_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1747_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1747_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1747_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1747_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1726 : std_logic_vector(31 downto 0);
    signal arrayidx81_1749 : std_logic_vector(31 downto 0);
    signal arrayidx81_1750_delayed_6_0_1752 : std_logic_vector(31 downto 0);
    signal call11_1519 : std_logic_vector(15 downto 0);
    signal call13_1522 : std_logic_vector(15 downto 0);
    signal call14_1525 : std_logic_vector(15 downto 0);
    signal call15_1528 : std_logic_vector(15 downto 0);
    signal call16_1541 : std_logic_vector(15 downto 0);
    signal call18_1553 : std_logic_vector(15 downto 0);
    signal call1_1504 : std_logic_vector(15 downto 0);
    signal call20_1556 : std_logic_vector(15 downto 0);
    signal call22_1559 : std_logic_vector(15 downto 0);
    signal call3_1507 : std_logic_vector(15 downto 0);
    signal call5_1510 : std_logic_vector(15 downto 0);
    signal call7_1513 : std_logic_vector(15 downto 0);
    signal call9_1516 : std_logic_vector(15 downto 0);
    signal call_1501 : std_logic_vector(15 downto 0);
    signal cmp104_1809 : std_logic_vector(0 downto 0);
    signal cmp116_1837 : std_logic_vector(0 downto 0);
    signal cmp_1770 : std_logic_vector(0 downto 0);
    signal conv111_1832 : std_logic_vector(31 downto 0);
    signal conv114_1606 : std_logic_vector(31 downto 0);
    signal conv17_1545 : std_logic_vector(31 downto 0);
    signal conv61_1687 : std_logic_vector(63 downto 0);
    signal conv64_1586 : std_logic_vector(63 downto 0);
    signal conv66_1691 : std_logic_vector(63 downto 0);
    signal conv69_1590 : std_logic_vector(63 downto 0);
    signal conv71_1695 : std_logic_vector(63 downto 0);
    signal conv90_1760 : std_logic_vector(31 downto 0);
    signal conv92_1602 : std_logic_vector(31 downto 0);
    signal conv_1532 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1790 : std_logic_vector(15 downto 0);
    signal idxprom80_1742 : std_logic_vector(63 downto 0);
    signal idxprom_1719 : std_logic_vector(63 downto 0);
    signal inc108_1813 : std_logic_vector(15 downto 0);
    signal inc108x_xinput_dim0x_x1_1821 : std_logic_vector(15 downto 0);
    signal inc_1796 : std_logic_vector(15 downto 0);
    signal indvar_1638 : std_logic_vector(31 downto 0);
    signal indvar_at_entry_1615 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1843 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1_1653 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_1804_delayed_3_0_1816 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_1630 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0_1804 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1648 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1790_delayed_2_0_1799 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_at_entry_1625 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1828 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0_1786 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1643 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_at_entry_1620 : std_logic_vector(15 downto 0);
    signal mul50_1678 : std_logic_vector(15 downto 0);
    signal mul72_1700 : std_logic_vector(63 downto 0);
    signal mul74_1710 : std_logic_vector(63 downto 0);
    signal mul_1668 : std_logic_vector(15 downto 0);
    signal ptr_deref_1729_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1729_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1729_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1729_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1729_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1754_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1754_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1754_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1754_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1754_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1754_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1538 : std_logic_vector(31 downto 0);
    signal shr115129_1612 : std_logic_vector(31 downto 0);
    signal shr_1736 : std_logic_vector(63 downto 0);
    signal sub44_1673 : std_logic_vector(15 downto 0);
    signal sub57_1582 : std_logic_vector(15 downto 0);
    signal sub58_1683 : std_logic_vector(15 downto 0);
    signal sub86_1596 : std_logic_vector(15 downto 0);
    signal sub_1571 : std_logic_vector(15 downto 0);
    signal tmp78_1730 : std_logic_vector(63 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1564_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1600_wire : std_logic_vector(31 downto 0);
    signal type_cast_1610_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1641_wire : std_logic_vector(31 downto 0);
    signal type_cast_1646_wire : std_logic_vector(15 downto 0);
    signal type_cast_1651_wire : std_logic_vector(15 downto 0);
    signal type_cast_1656_wire : std_logic_vector(15 downto 0);
    signal type_cast_1734_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1740_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1762_1762_delayed_2_0_1764 : std_logic_vector(31 downto 0);
    signal type_cast_1767_wire : std_logic_vector(31 downto 0);
    signal type_cast_1774_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1784_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1794_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1825_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1841_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1858_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_whilex_xend_taken_1846 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_1724_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1724_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1724_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1724_resized_base_address <= "00000000000000";
    array_obj_ref_1747_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1747_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1747_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1747_resized_base_address <= "00000000000000";
    indvar_at_entry_1615 <= "00000000000000000000000000000000";
    input_dim0x_x1_at_entry_1630 <= "0000000000000000";
    input_dim1x_x1_at_entry_1625 <= "0000000000000000";
    input_dim2x_x1_at_entry_1620 <= "0000000000000000";
    ptr_deref_1729_word_offset_0 <= "00000000000000";
    ptr_deref_1754_word_offset_0 <= "00000000000000";
    type_cast_1536_wire_constant <= "00000000000000000000000000010000";
    type_cast_1564_wire_constant <= "1111111111111111";
    type_cast_1575_wire_constant <= "1111111111111111";
    type_cast_1594_wire_constant <= "1111111111111100";
    type_cast_1610_wire_constant <= "00000000000000000000000000000010";
    type_cast_1734_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1740_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1774_wire_constant <= "0000000000000100";
    type_cast_1784_wire_constant <= "0000000000000000";
    type_cast_1794_wire_constant <= "0000000000000001";
    type_cast_1825_wire_constant <= "0000000000000000";
    type_cast_1841_wire_constant <= "00000000000000000000000000000001";
    type_cast_1858_wire_constant <= "0000000000000001";
    phi_stmt_1638: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1641_wire & indvar_at_entry_1615;
      req <= phi_stmt_1638_req_0 & phi_stmt_1638_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1638",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1638_ack_0,
          idata => idata,
          odata => indvar_1638,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1638
    phi_stmt_1643: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1646_wire & input_dim2x_x1_at_entry_1620;
      req <= phi_stmt_1643_req_0 & phi_stmt_1643_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1643",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1643_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1643,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1643
    phi_stmt_1648: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1651_wire & input_dim1x_x1_at_entry_1625;
      req <= phi_stmt_1648_req_0 & phi_stmt_1648_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1648",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1648_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1648,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1648
    phi_stmt_1653: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1656_wire & input_dim0x_x1_at_entry_1630;
      req <= phi_stmt_1653_req_0 & phi_stmt_1653_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1653",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1653_ack_0,
          idata => idata,
          odata => input_dim0x_x1_1653,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1653
    -- flow-through select operator MUX_1785_inst
    input_dim2x_x0_1786 <= add96_1773_delayed_1_0_1779 when (cmp_1770(0) /=  '0') else type_cast_1784_wire_constant;
    -- flow-through select operator MUX_1827_inst
    input_dim1x_x2_1828 <= type_cast_1825_wire_constant when (cmp104_1809(0) /=  '0') else input_dim1x_x0_1804;
    W_add96_1773_delayed_1_0_1777_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add96_1773_delayed_1_0_1777_inst_req_0;
      W_add96_1773_delayed_1_0_1777_inst_ack_0<= wack(0);
      rreq(0) <= W_add96_1773_delayed_1_0_1777_inst_req_1;
      W_add96_1773_delayed_1_0_1777_inst_ack_1<= rack(0);
      W_add96_1773_delayed_1_0_1777_inst : InterlockBuffer generic map ( -- 
        name => "W_add96_1773_delayed_1_0_1777_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add96_1776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add96_1773_delayed_1_0_1779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx81_1750_delayed_6_0_1750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx81_1750_delayed_6_0_1750_inst_req_0;
      W_arrayidx81_1750_delayed_6_0_1750_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx81_1750_delayed_6_0_1750_inst_req_1;
      W_arrayidx81_1750_delayed_6_0_1750_inst_ack_1<= rack(0);
      W_arrayidx81_1750_delayed_6_0_1750_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx81_1750_delayed_6_0_1750_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx81_1749,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx81_1750_delayed_6_0_1752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim0x_x1_1804_delayed_3_0_1814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim0x_x1_1804_delayed_3_0_1814_inst_req_0;
      W_input_dim0x_x1_1804_delayed_3_0_1814_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim0x_x1_1804_delayed_3_0_1814_inst_req_1;
      W_input_dim0x_x1_1804_delayed_3_0_1814_inst_ack_1<= rack(0);
      W_input_dim0x_x1_1804_delayed_3_0_1814_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim0x_x1_1804_delayed_3_0_1814_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_1653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_1804_delayed_3_0_1816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim1x_x1_1790_delayed_2_0_1797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim1x_x1_1790_delayed_2_0_1797_inst_req_0;
      W_input_dim1x_x1_1790_delayed_2_0_1797_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim1x_x1_1790_delayed_2_0_1797_inst_req_1;
      W_input_dim1x_x1_1790_delayed_2_0_1797_inst_ack_1<= rack(0);
      W_input_dim1x_x1_1790_delayed_2_0_1797_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim1x_x1_1790_delayed_2_0_1797_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim1x_x1_1790_delayed_2_0_1799,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_1844_inst
    process(cmp116_1837) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp116_1837(0 downto 0);
      whilex_xbody_whilex_xend_taken_1846 <= tmp_var; -- 
    end process;
    addr_of_1725_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1725_final_reg_req_0;
      addr_of_1725_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1725_final_reg_req_1;
      addr_of_1725_final_reg_ack_1<= rack(0);
      addr_of_1725_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1725_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1724_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1726,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1748_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1748_final_reg_req_0;
      addr_of_1748_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1748_final_reg_req_1;
      addr_of_1748_final_reg_ack_1<= rack(0);
      addr_of_1748_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1748_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1747_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx81_1749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1531_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1531_inst_req_0;
      type_cast_1531_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1531_inst_req_1;
      type_cast_1531_inst_ack_1<= rack(0);
      type_cast_1531_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1531_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1528,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1544_inst_req_0;
      type_cast_1544_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1544_inst_req_1;
      type_cast_1544_inst_ack_1<= rack(0);
      type_cast_1544_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1544_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1585_inst_req_0;
      type_cast_1585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1585_inst_req_1;
      type_cast_1585_inst_ack_1<= rack(0);
      type_cast_1585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1559,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1589_inst_req_0;
      type_cast_1589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1589_inst_req_1;
      type_cast_1589_inst_ack_1<= rack(0);
      type_cast_1589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1601_inst_req_0;
      type_cast_1601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1601_inst_req_1;
      type_cast_1601_inst_ack_1<= rack(0);
      type_cast_1601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1600_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv92_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1605_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1605_inst_req_0;
      type_cast_1605_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1605_inst_req_1;
      type_cast_1605_inst_ack_1<= rack(0);
      type_cast_1605_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1605_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv114_1606,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1641_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1641_inst_req_0;
      type_cast_1641_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1641_inst_req_1;
      type_cast_1641_inst_ack_1<= rack(0);
      type_cast_1641_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1641_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1843,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1641_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1646_inst_req_0;
      type_cast_1646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1646_inst_req_1;
      type_cast_1646_inst_ack_1<= rack(0);
      type_cast_1646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1646_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0_1786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1646_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1651_inst_req_0;
      type_cast_1651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1651_inst_req_1;
      type_cast_1651_inst_ack_1<= rack(0);
      type_cast_1651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1651_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1651_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1656_inst_req_0;
      type_cast_1656_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1656_inst_req_1;
      type_cast_1656_inst_ack_1<= rack(0);
      type_cast_1656_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1656_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc108x_xinput_dim0x_x1_1821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1656_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1686_inst_req_0;
      type_cast_1686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1686_inst_req_1;
      type_cast_1686_inst_ack_1<= rack(0);
      type_cast_1686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1643,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1690_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1690_inst_req_0;
      type_cast_1690_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1690_inst_req_1;
      type_cast_1690_inst_ack_1<= rack(0);
      type_cast_1690_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1690_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1691,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1694_inst_req_0;
      type_cast_1694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1694_inst_req_1;
      type_cast_1694_inst_ack_1<= rack(0);
      type_cast_1694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1718_inst_req_0;
      type_cast_1718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1718_inst_req_1;
      type_cast_1718_inst_ack_1<= rack(0);
      type_cast_1718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_src_0x_x0_1663,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1759_inst_req_0;
      type_cast_1759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1759_inst_req_1;
      type_cast_1759_inst_ack_1<= rack(0);
      type_cast_1759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1759_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1643,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1763_inst_req_0;
      type_cast_1763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1763_inst_req_1;
      type_cast_1763_inst_ack_1<= rack(0);
      type_cast_1763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1763_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv92_1602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1762_1762_delayed_2_0_1764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1767_inst
    process(conv90_1760) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv90_1760(31 downto 0);
      type_cast_1767_wire <= tmp_var; -- 
    end process;
    type_cast_1789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1789_inst_req_0;
      type_cast_1789_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1789_inst_req_1;
      type_cast_1789_inst_ack_1<= rack(0);
      type_cast_1789_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1789_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_1770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_18_1790,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1812_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1812_inst_req_0;
      type_cast_1812_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1812_inst_req_1;
      type_cast_1812_inst_ack_1<= rack(0);
      type_cast_1812_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1812_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp104_1809,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc108_1813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1831_inst_req_0;
      type_cast_1831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1831_inst_req_1;
      type_cast_1831_inst_ack_1<= rack(0);
      type_cast_1831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc108x_xinput_dim0x_x1_1821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1724_index_1_rename
    process(R_idxprom_1723_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1723_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1723_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1724_index_1_resize
    process(idxprom_1719) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1719;
      ov := iv(13 downto 0);
      R_idxprom_1723_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1724_root_address_inst
    process(array_obj_ref_1724_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1724_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1724_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1747_index_1_rename
    process(R_idxprom80_1746_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom80_1746_resized;
      ov(13 downto 0) := iv;
      R_idxprom80_1746_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1747_index_1_resize
    process(idxprom80_1742) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom80_1742;
      ov := iv(13 downto 0);
      R_idxprom80_1746_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1747_root_address_inst
    process(array_obj_ref_1747_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1747_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1747_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1729_addr_0
    process(ptr_deref_1729_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1729_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1729_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1729_base_resize
    process(arrayidx77_1726) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1726;
      ov := iv(13 downto 0);
      ptr_deref_1729_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1729_gather_scatter
    process(ptr_deref_1729_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1729_data_0;
      ov(63 downto 0) := iv;
      tmp78_1730 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1729_root_address_inst
    process(ptr_deref_1729_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1729_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1729_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1754_addr_0
    process(ptr_deref_1754_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1754_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1754_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1754_base_resize
    process(arrayidx81_1750_delayed_6_0_1752) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx81_1750_delayed_6_0_1752;
      ov := iv(13 downto 0);
      ptr_deref_1754_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1754_gather_scatter
    process(tmp78_1730) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1730;
      ov(63 downto 0) := iv;
      ptr_deref_1754_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1754_root_address_inst
    process(ptr_deref_1754_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1754_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1754_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_1636_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1849_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1636_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1636_branch_req_0,
          ack0 => do_while_stmt_1636_branch_ack_0,
          ack1 => do_while_stmt_1636_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1850_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_1846;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1850_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1850_branch_req_0,
          ack0 => if_stmt_1850_branch_ack_0,
          ack1 => if_stmt_1850_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1565_inst
    process(call7_1513) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1513, type_cast_1564_wire_constant, tmp_var);
      add41_1566 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1576_inst
    process(call9_1516) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1516, type_cast_1575_wire_constant, tmp_var);
      add54_1577 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1595_inst
    process(call3_1507) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call3_1507, type_cast_1594_wire_constant, tmp_var);
      sub86_1596 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1672_inst
    process(sub_1571, mul_1668) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1571, mul_1668, tmp_var);
      sub44_1673 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1682_inst
    process(sub57_1582, mul50_1678) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1582, mul50_1678, tmp_var);
      sub58_1683 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1775_inst
    process(input_dim2x_x1_1643) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1643, type_cast_1774_wire_constant, tmp_var);
      add96_1776 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1803_inst
    process(inc_1796, input_dim1x_x1_1790_delayed_2_0_1799) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc_1796, input_dim1x_x1_1790_delayed_2_0_1799, tmp_var);
      input_dim1x_x0_1804 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1820_inst
    process(inc108_1813, input_dim0x_x1_1804_delayed_3_0_1816) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc108_1813, input_dim0x_x1_1804_delayed_3_0_1816, tmp_var);
      inc108x_xinput_dim0x_x1_1821 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1662_inst
    process(add_1550, indvar_1638) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1550, indvar_1638, tmp_var);
      add_src_0x_x0_1663 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1842_inst
    process(indvar_1638) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1638, type_cast_1841_wire_constant, tmp_var);
      indvarx_xnext_1843 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1704_inst
    process(mul72_1700, conv66_1691) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1700, conv66_1691, tmp_var);
      add73_1705 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1714_inst
    process(mul74_1710, conv61_1687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1710, conv61_1687, tmp_var);
      add75_1715 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1741_inst
    process(shr_1736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr_1736, type_cast_1740_wire_constant, tmp_var);
      idxprom80_1742 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1808_inst
    process(input_dim1x_x0_1804, call1_1504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1x_x0_1804, call1_1504, tmp_var);
      cmp104_1809 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1836_inst
    process(conv111_1832, shr115129_1612) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv111_1832, shr115129_1612, tmp_var);
      cmp116_1837 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1611_inst
    process(conv114_1606) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv114_1606, type_cast_1610_wire_constant, tmp_var);
      shr115129_1612 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1735_inst
    process(add75_1715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1715, type_cast_1734_wire_constant, tmp_var);
      shr_1736 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1667_inst
    process(input_dim0x_x1_1653, call13_1522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x1_1653, call13_1522, tmp_var);
      mul_1668 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1677_inst
    process(input_dim1x_x1_1648, call13_1522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1648, call13_1522, tmp_var);
      mul50_1678 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1699_inst
    process(conv71_1695, conv69_1590) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1695, conv69_1590, tmp_var);
      mul72_1700 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1709_inst
    process(add73_1705, conv64_1586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1705, conv64_1586, tmp_var);
      mul74_1710 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1849_inst
    process(cmp116_1837) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp116_1837, tmp_var);
      NOT_u1_u1_1849_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u32_u32_1549_inst
    process(shl_1538, conv17_1545) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1538, conv17_1545, tmp_var);
      add_1550 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1537_inst
    process(conv_1532) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1532, type_cast_1536_wire_constant, tmp_var);
      shl_1538 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1769_inst
    process(type_cast_1767_wire, type_cast_1762_1762_delayed_2_0_1764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1767_wire, type_cast_1762_1762_delayed_2_0_1764, tmp_var);
      cmp_1770 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1570_inst
    process(add41_1566, call14_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1566, call14_1525, tmp_var);
      sub_1571 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1581_inst
    process(add54_1577, call14_1525) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1577, call14_1525, tmp_var);
      sub57_1582 <= tmp_var; --
    end process;
    -- binary operator XOR_u16_u16_1795_inst
    process(iNsTr_18_1790) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntXor_proc(iNsTr_18_1790, type_cast_1794_wire_constant, tmp_var);
      inc_1796 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1724_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1723_scaled;
      array_obj_ref_1724_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1724_index_offset_req_0;
      array_obj_ref_1724_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1724_index_offset_req_1;
      array_obj_ref_1724_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1747_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom80_1746_scaled;
      array_obj_ref_1747_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1747_index_offset_req_0;
      array_obj_ref_1747_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1747_index_offset_req_1;
      array_obj_ref_1747_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- unary operator type_cast_1600_inst
    process(sub86_1596) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", sub86_1596, tmp_var);
      type_cast_1600_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1729_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1729_load_0_req_0;
      ptr_deref_1729_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1729_load_0_req_1;
      ptr_deref_1729_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1729_word_address_0;
      ptr_deref_1729_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1754_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1754_store_0_req_0;
      ptr_deref_1754_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1754_store_0_req_1;
      ptr_deref_1754_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1754_word_address_0;
      data_in <= ptr_deref_1754_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1500_inst RPIPE_Block0_start_1503_inst RPIPE_Block0_start_1506_inst RPIPE_Block0_start_1509_inst RPIPE_Block0_start_1512_inst RPIPE_Block0_start_1515_inst RPIPE_Block0_start_1518_inst RPIPE_Block0_start_1521_inst RPIPE_Block0_start_1524_inst RPIPE_Block0_start_1527_inst RPIPE_Block0_start_1540_inst RPIPE_Block0_start_1552_inst RPIPE_Block0_start_1555_inst RPIPE_Block0_start_1558_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1500_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1503_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1506_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1509_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1512_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1515_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1518_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1521_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1524_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1527_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1540_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1552_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1555_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1558_inst_req_0;
      RPIPE_Block0_start_1500_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1503_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1506_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1509_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1512_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1515_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1518_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1521_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1524_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1527_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1540_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1552_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1555_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1558_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1500_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1503_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1506_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1509_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1512_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1515_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1518_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1521_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1524_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1527_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1540_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1552_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1555_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1558_inst_req_1;
      RPIPE_Block0_start_1500_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1503_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1506_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1509_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1512_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1515_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1518_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1521_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1524_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1527_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1540_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1552_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1555_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1558_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_1501 <= data_out(223 downto 208);
      call1_1504 <= data_out(207 downto 192);
      call3_1507 <= data_out(191 downto 176);
      call5_1510 <= data_out(175 downto 160);
      call7_1513 <= data_out(159 downto 144);
      call9_1516 <= data_out(143 downto 128);
      call11_1519 <= data_out(127 downto 112);
      call13_1522 <= data_out(111 downto 96);
      call14_1525 <= data_out(95 downto 80);
      call15_1528 <= data_out(79 downto 64);
      call16_1541 <= data_out(63 downto 48);
      call18_1553 <= data_out(47 downto 32);
      call20_1556 <= data_out(31 downto 16);
      call22_1559 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1856_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1856_inst_req_0;
      WPIPE_Block0_done_1856_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1856_inst_req_1;
      WPIPE_Block0_done_1856_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1858_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4715_start: Boolean;
  signal convTransposeB_CP_4715_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2018_inst_req_1 : boolean;
  signal ptr_deref_2100_load_0_ack_1 : boolean;
  signal W_arrayidx86_2106_delayed_6_0_2121_inst_req_0 : boolean;
  signal type_cast_2023_inst_ack_1 : boolean;
  signal type_cast_2057_inst_req_0 : boolean;
  signal type_cast_2018_inst_ack_0 : boolean;
  signal type_cast_2018_inst_req_0 : boolean;
  signal ptr_deref_2100_load_0_req_1 : boolean;
  signal type_cast_2089_inst_ack_1 : boolean;
  signal addr_of_2096_final_reg_ack_1 : boolean;
  signal input_dim0x_x1_at_entry_2002_2028_buf_ack_1 : boolean;
  signal input_dim0x_x1_at_entry_2002_2028_buf_req_1 : boolean;
  signal input_dim0x_x1_at_entry_2002_2028_buf_ack_0 : boolean;
  signal input_dim0x_x1_at_entry_2002_2028_buf_req_0 : boolean;
  signal type_cast_2089_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1867_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_req_1 : boolean;
  signal addr_of_2096_final_reg_req_0 : boolean;
  signal addr_of_2096_final_reg_ack_0 : boolean;
  signal RPIPE_Block1_start_1867_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1867_inst_req_0 : boolean;
  signal type_cast_2023_inst_req_1 : boolean;
  signal ptr_deref_2125_store_0_req_0 : boolean;
  signal RPIPE_Block1_start_1873_inst_ack_1 : boolean;
  signal type_cast_2089_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1873_inst_req_0 : boolean;
  signal type_cast_2018_inst_ack_1 : boolean;
  signal addr_of_2119_final_reg_ack_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1879_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1879_inst_req_0 : boolean;
  signal type_cast_2089_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1870_inst_req_0 : boolean;
  signal addr_of_2119_final_reg_req_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_ack_0 : boolean;
  signal type_cast_2023_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1879_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1879_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1876_inst_ack_1 : boolean;
  signal addr_of_2119_final_reg_req_0 : boolean;
  signal RPIPE_Block1_start_1882_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1882_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1882_inst_ack_0 : boolean;
  signal type_cast_2023_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1882_inst_req_0 : boolean;
  signal type_cast_2057_inst_req_1 : boolean;
  signal ptr_deref_2125_store_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1885_inst_req_0 : boolean;
  signal type_cast_2057_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1885_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1885_inst_ack_1 : boolean;
  signal type_cast_2130_inst_req_0 : boolean;
  signal type_cast_2130_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1885_inst_ack_0 : boolean;
  signal type_cast_2130_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_req_0 : boolean;
  signal addr_of_2119_final_reg_ack_0 : boolean;
  signal addr_of_2096_final_reg_req_1 : boolean;
  signal type_cast_2130_inst_ack_1 : boolean;
  signal W_arrayidx86_2106_delayed_6_0_2121_inst_ack_0 : boolean;
  signal ptr_deref_2125_store_0_ack_1 : boolean;
  signal array_obj_ref_2095_index_offset_ack_1 : boolean;
  signal RPIPE_Block1_start_1888_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1888_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1888_inst_req_1 : boolean;
  signal type_cast_2065_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1888_inst_ack_1 : boolean;
  signal ptr_deref_2125_store_0_req_1 : boolean;
  signal type_cast_2027_inst_ack_1 : boolean;
  signal array_obj_ref_2095_index_offset_req_1 : boolean;
  signal type_cast_2027_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1891_inst_req_0 : boolean;
  signal type_cast_2065_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1891_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1891_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1891_inst_ack_1 : boolean;
  signal array_obj_ref_2118_index_offset_ack_1 : boolean;
  signal array_obj_ref_2118_index_offset_req_1 : boolean;
  signal RPIPE_Block1_start_1894_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1894_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1894_inst_req_1 : boolean;
  signal type_cast_2065_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1894_inst_ack_1 : boolean;
  signal array_obj_ref_2118_index_offset_ack_0 : boolean;
  signal array_obj_ref_2118_index_offset_req_0 : boolean;
  signal type_cast_2027_inst_ack_0 : boolean;
  signal array_obj_ref_2095_index_offset_ack_0 : boolean;
  signal type_cast_2027_inst_req_0 : boolean;
  signal type_cast_1898_inst_req_0 : boolean;
  signal type_cast_2065_inst_req_0 : boolean;
  signal type_cast_1898_inst_ack_0 : boolean;
  signal type_cast_1898_inst_req_1 : boolean;
  signal type_cast_1898_inst_ack_1 : boolean;
  signal phi_stmt_2019_ack_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1907_inst_ack_1 : boolean;
  signal phi_stmt_2019_req_0 : boolean;
  signal phi_stmt_2019_req_1 : boolean;
  signal array_obj_ref_2095_index_offset_req_0 : boolean;
  signal type_cast_1911_inst_req_0 : boolean;
  signal type_cast_1911_inst_ack_0 : boolean;
  signal type_cast_1911_inst_req_1 : boolean;
  signal type_cast_1911_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1919_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1919_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1919_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1919_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1922_inst_req_0 : boolean;
  signal type_cast_2061_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1922_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1922_inst_req_1 : boolean;
  signal type_cast_2061_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1922_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1925_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1925_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1925_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1925_inst_ack_1 : boolean;
  signal type_cast_1958_inst_req_0 : boolean;
  signal type_cast_2061_inst_ack_0 : boolean;
  signal type_cast_1958_inst_ack_0 : boolean;
  signal ptr_deref_2100_load_0_ack_0 : boolean;
  signal ptr_deref_2100_load_0_req_0 : boolean;
  signal type_cast_1958_inst_req_1 : boolean;
  signal type_cast_2061_inst_req_0 : boolean;
  signal type_cast_1958_inst_ack_1 : boolean;
  signal type_cast_1962_inst_req_0 : boolean;
  signal type_cast_1962_inst_ack_0 : boolean;
  signal type_cast_1962_inst_req_1 : boolean;
  signal type_cast_1962_inst_ack_1 : boolean;
  signal type_cast_1973_inst_req_0 : boolean;
  signal type_cast_1973_inst_ack_0 : boolean;
  signal type_cast_1973_inst_req_1 : boolean;
  signal type_cast_1973_inst_ack_1 : boolean;
  signal W_arrayidx86_2106_delayed_6_0_2121_inst_ack_1 : boolean;
  signal W_arrayidx86_2106_delayed_6_0_2121_inst_req_1 : boolean;
  signal type_cast_1977_inst_req_0 : boolean;
  signal type_cast_1977_inst_ack_0 : boolean;
  signal type_cast_1977_inst_req_1 : boolean;
  signal type_cast_1977_inst_ack_1 : boolean;
  signal phi_stmt_2024_ack_0 : boolean;
  signal do_while_stmt_2007_branch_req_0 : boolean;
  signal type_cast_2057_inst_ack_1 : boolean;
  signal phi_stmt_2024_req_1 : boolean;
  signal phi_stmt_2024_req_0 : boolean;
  signal phi_stmt_2009_req_0 : boolean;
  signal phi_stmt_2009_req_1 : boolean;
  signal phi_stmt_2009_ack_0 : boolean;
  signal type_cast_2012_inst_req_0 : boolean;
  signal type_cast_2012_inst_ack_0 : boolean;
  signal type_cast_2012_inst_req_1 : boolean;
  signal type_cast_2012_inst_ack_1 : boolean;
  signal phi_stmt_2014_req_1 : boolean;
  signal phi_stmt_2014_req_0 : boolean;
  signal phi_stmt_2014_ack_0 : boolean;
  signal type_cast_2134_inst_req_0 : boolean;
  signal type_cast_2134_inst_ack_0 : boolean;
  signal type_cast_2134_inst_req_1 : boolean;
  signal type_cast_2134_inst_ack_1 : boolean;
  signal W_add101_2129_delayed_1_0_2148_inst_req_0 : boolean;
  signal W_add101_2129_delayed_1_0_2148_inst_ack_0 : boolean;
  signal W_add101_2129_delayed_1_0_2148_inst_req_1 : boolean;
  signal W_add101_2129_delayed_1_0_2148_inst_ack_1 : boolean;
  signal type_cast_2160_inst_req_0 : boolean;
  signal type_cast_2160_inst_ack_0 : boolean;
  signal type_cast_2160_inst_req_1 : boolean;
  signal type_cast_2160_inst_ack_1 : boolean;
  signal W_input_dim1x_x1_2146_delayed_2_0_2168_inst_req_0 : boolean;
  signal W_input_dim1x_x1_2146_delayed_2_0_2168_inst_ack_0 : boolean;
  signal W_input_dim1x_x1_2146_delayed_2_0_2168_inst_req_1 : boolean;
  signal W_input_dim1x_x1_2146_delayed_2_0_2168_inst_ack_1 : boolean;
  signal type_cast_2183_inst_req_0 : boolean;
  signal type_cast_2183_inst_ack_0 : boolean;
  signal type_cast_2183_inst_req_1 : boolean;
  signal type_cast_2183_inst_ack_1 : boolean;
  signal W_input_dim0x_x1_2160_delayed_3_0_2185_inst_req_0 : boolean;
  signal W_input_dim0x_x1_2160_delayed_3_0_2185_inst_ack_0 : boolean;
  signal W_input_dim0x_x1_2160_delayed_3_0_2185_inst_req_1 : boolean;
  signal W_input_dim0x_x1_2160_delayed_3_0_2185_inst_ack_1 : boolean;
  signal type_cast_2202_inst_req_0 : boolean;
  signal type_cast_2202_inst_ack_0 : boolean;
  signal type_cast_2202_inst_req_1 : boolean;
  signal type_cast_2202_inst_ack_1 : boolean;
  signal do_while_stmt_2007_branch_ack_0 : boolean;
  signal do_while_stmt_2007_branch_ack_1 : boolean;
  signal if_stmt_2221_branch_req_0 : boolean;
  signal if_stmt_2221_branch_ack_1 : boolean;
  signal if_stmt_2221_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2227_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2227_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2227_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2227_inst_ack_1 : boolean;
  signal type_cast_2005_inst_req_0 : boolean;
  signal type_cast_2005_inst_ack_0 : boolean;
  signal type_cast_2005_inst_req_1 : boolean;
  signal type_cast_2005_inst_ack_1 : boolean;
  signal phi_stmt_2002_req_0 : boolean;
  signal phi_stmt_2002_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4715_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4715_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4715_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4715_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4715: Block -- control-path 
    signal convTransposeB_CP_4715_elements: BooleanArray(226 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4715_elements(0) <= convTransposeB_CP_4715_start;
    convTransposeB_CP_4715_symbol <= convTransposeB_CP_4715_elements(222);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1865/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926__entry__
      -- CP-element group 0: 	 branch_block_stmt_1865/branch_block_stmt_1865__entry__
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/$entry
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Update/cr
      -- 
    rr_4749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(0), ack => RPIPE_Block1_start_1867_inst_req_0); -- 
    cr_4894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(0), ack => type_cast_1898_inst_req_1); -- 
    cr_4922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(0), ack => type_cast_1911_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	218 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	219 
    -- CP-element group 1: 	220 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221__entry__
      -- CP-element group 1: 	 branch_block_stmt_1865/do_while_stmt_2007__exit__
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1865/R_whilex_xbody_whilex_xend_taken_2222_place
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1865/if_stmt_2221_else_link/$entry
      -- 
    branch_req_5622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(1), ack => if_stmt_2221_branch_req_0); -- 
    convTransposeB_CP_4715_elements(1) <= convTransposeB_CP_4715_elements(218);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_sample_completed_
      -- 
    ra_4750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1867_inst_ack_0, ack => convTransposeB_CP_4715_elements(2)); -- 
    cr_4754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(2), ack => RPIPE_Block1_start_1867_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1867_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_sample_start_
      -- 
    ca_4755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1867_inst_ack_1, ack => convTransposeB_CP_4715_elements(3)); -- 
    rr_4763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(3), ack => RPIPE_Block1_start_1870_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_sample_completed_
      -- 
    ra_4764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1870_inst_ack_0, ack => convTransposeB_CP_4715_elements(4)); -- 
    cr_4768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(4), ack => RPIPE_Block1_start_1870_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1870_update_completed_
      -- 
    ca_4769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1870_inst_ack_1, ack => convTransposeB_CP_4715_elements(5)); -- 
    rr_4777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(5), ack => RPIPE_Block1_start_1873_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_sample_completed_
      -- 
    ra_4778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1873_inst_ack_0, ack => convTransposeB_CP_4715_elements(6)); -- 
    cr_4782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(6), ack => RPIPE_Block1_start_1873_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1873_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Sample/rr
      -- 
    ca_4783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1873_inst_ack_1, ack => convTransposeB_CP_4715_elements(7)); -- 
    rr_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(7), ack => RPIPE_Block1_start_1876_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Update/$entry
      -- 
    ra_4792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1876_inst_ack_0, ack => convTransposeB_CP_4715_elements(8)); -- 
    cr_4796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(8), ack => RPIPE_Block1_start_1876_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1876_Update/$exit
      -- 
    ca_4797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1876_inst_ack_1, ack => convTransposeB_CP_4715_elements(9)); -- 
    rr_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(9), ack => RPIPE_Block1_start_1879_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_sample_completed_
      -- 
    ra_4806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1879_inst_ack_0, ack => convTransposeB_CP_4715_elements(10)); -- 
    cr_4810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(10), ack => RPIPE_Block1_start_1879_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1879_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_sample_start_
      -- 
    ca_4811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1879_inst_ack_1, ack => convTransposeB_CP_4715_elements(11)); -- 
    rr_4819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(11), ack => RPIPE_Block1_start_1882_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_sample_completed_
      -- 
    ra_4820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1882_inst_ack_0, ack => convTransposeB_CP_4715_elements(12)); -- 
    cr_4824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(12), ack => RPIPE_Block1_start_1882_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1882_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Sample/$entry
      -- 
    ca_4825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1882_inst_ack_1, ack => convTransposeB_CP_4715_elements(13)); -- 
    rr_4833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(13), ack => RPIPE_Block1_start_1885_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_update_start_
      -- 
    ra_4834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1885_inst_ack_0, ack => convTransposeB_CP_4715_elements(14)); -- 
    cr_4838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(14), ack => RPIPE_Block1_start_1885_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1885_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Sample/rr
      -- 
    ca_4839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1885_inst_ack_1, ack => convTransposeB_CP_4715_elements(15)); -- 
    rr_4847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(15), ack => RPIPE_Block1_start_1888_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Update/cr
      -- 
    ra_4848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1888_inst_ack_0, ack => convTransposeB_CP_4715_elements(16)); -- 
    cr_4852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(16), ack => RPIPE_Block1_start_1888_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1888_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Sample/rr
      -- 
    ca_4853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1888_inst_ack_1, ack => convTransposeB_CP_4715_elements(17)); -- 
    rr_4861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(17), ack => RPIPE_Block1_start_1891_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Update/cr
      -- 
    ra_4862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1891_inst_ack_0, ack => convTransposeB_CP_4715_elements(18)); -- 
    cr_4866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(18), ack => RPIPE_Block1_start_1891_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1891_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Sample/rr
      -- 
    ca_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1891_inst_ack_1, ack => convTransposeB_CP_4715_elements(19)); -- 
    rr_4875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(19), ack => RPIPE_Block1_start_1894_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Update/cr
      -- 
    ra_4876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1894_inst_ack_0, ack => convTransposeB_CP_4715_elements(20)); -- 
    cr_4880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(20), ack => RPIPE_Block1_start_1894_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1894_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Sample/rr
      -- 
    ca_4881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1894_inst_ack_1, ack => convTransposeB_CP_4715_elements(21)); -- 
    rr_4903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(21), ack => RPIPE_Block1_start_1907_inst_req_0); -- 
    rr_4889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(21), ack => type_cast_1898_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Sample/ra
      -- 
    ra_4890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1898_inst_ack_0, ack => convTransposeB_CP_4715_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1898_Update/ca
      -- 
    ca_4895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1898_inst_ack_1, ack => convTransposeB_CP_4715_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Update/cr
      -- 
    ra_4904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1907_inst_ack_0, ack => convTransposeB_CP_4715_elements(24)); -- 
    cr_4908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(24), ack => RPIPE_Block1_start_1907_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1907_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Sample/rr
      -- 
    ca_4909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1907_inst_ack_1, ack => convTransposeB_CP_4715_elements(25)); -- 
    rr_4917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(25), ack => type_cast_1911_inst_req_0); -- 
    rr_4931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(25), ack => RPIPE_Block1_start_1919_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Sample/ra
      -- 
    ra_4918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1911_inst_ack_0, ack => convTransposeB_CP_4715_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/type_cast_1911_Update/ca
      -- 
    ca_4923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1911_inst_ack_1, ack => convTransposeB_CP_4715_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Update/cr
      -- 
    ra_4932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1919_inst_ack_0, ack => convTransposeB_CP_4715_elements(28)); -- 
    cr_4936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(28), ack => RPIPE_Block1_start_1919_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1919_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Sample/rr
      -- 
    ca_4937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1919_inst_ack_1, ack => convTransposeB_CP_4715_elements(29)); -- 
    rr_4945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(29), ack => RPIPE_Block1_start_1922_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Update/cr
      -- 
    ra_4946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1922_inst_ack_0, ack => convTransposeB_CP_4715_elements(30)); -- 
    cr_4950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(30), ack => RPIPE_Block1_start_1922_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1922_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Sample/rr
      -- 
    ca_4951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1922_inst_ack_1, ack => convTransposeB_CP_4715_elements(31)); -- 
    rr_4959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(31), ack => RPIPE_Block1_start_1925_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Update/cr
      -- 
    ra_4960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1925_inst_ack_0, ack => convTransposeB_CP_4715_elements(32)); -- 
    cr_4964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(32), ack => RPIPE_Block1_start_1925_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/RPIPE_Block1_start_1925_Update/ca
      -- 
    ca_4965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1925_inst_ack_1, ack => convTransposeB_CP_4715_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984__entry__
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926__exit__
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1868_to_assign_stmt_1926/$exit
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Update/cr
      -- 
    rr_4976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1958_inst_req_0); -- 
    cr_4981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1958_inst_req_1); -- 
    rr_4990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1962_inst_req_0); -- 
    cr_4995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1962_inst_req_1); -- 
    rr_5004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1973_inst_req_0); -- 
    cr_5009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1973_inst_req_1); -- 
    rr_5018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1977_inst_req_0); -- 
    cr_5023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(34), ack => type_cast_1977_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(23) & convTransposeB_CP_4715_elements(27) & convTransposeB_CP_4715_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Sample/ra
      -- 
    ra_4977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1958_inst_ack_0, ack => convTransposeB_CP_4715_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1958_Update/ca
      -- 
    ca_4982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1958_inst_ack_1, ack => convTransposeB_CP_4715_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Sample/ra
      -- 
    ra_4991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1962_inst_ack_0, ack => convTransposeB_CP_4715_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1962_Update/ca
      -- 
    ca_4996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1962_inst_ack_1, ack => convTransposeB_CP_4715_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Sample/ra
      -- 
    ra_5005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1973_inst_ack_0, ack => convTransposeB_CP_4715_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1973_Update/ca
      -- 
    ca_5010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1973_inst_ack_1, ack => convTransposeB_CP_4715_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Sample/ra
      -- 
    ra_5019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1977_inst_ack_0, ack => convTransposeB_CP_4715_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/type_cast_1977_Update/ca
      -- 
    ca_5024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1977_inst_ack_1, ack => convTransposeB_CP_4715_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	223 
    -- CP-element group 43: 	224 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984__exit__
      -- CP-element group 43: 	 branch_block_stmt_1865/assign_stmt_1933_to_assign_stmt_1984/$exit
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Update/cr
      -- 
    rr_5668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(43), ack => type_cast_2005_inst_req_0); -- 
    cr_5673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(43), ack => type_cast_2005_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(36) & convTransposeB_CP_4715_elements(38) & convTransposeB_CP_4715_elements(40) & convTransposeB_CP_4715_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	226 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1865/do_while_stmt_2007/$entry
      -- CP-element group 44: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007__entry__
      -- 
    convTransposeB_CP_4715_elements(44) <= convTransposeB_CP_4715_elements(226);
    -- CP-element group 45:  merge  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	218 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007__exit__
      -- 
    -- Element group convTransposeB_CP_4715_elements(45) is bound as output of CP function.
    -- CP-element group 46:  merge  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_back
      -- 
    -- Element group convTransposeB_CP_4715_elements(46) is bound as output of CP function.
    -- CP-element group 47:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	52 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	217 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1865/do_while_stmt_2007/condition_done
      -- CP-element group 47: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_exit/$entry
      -- CP-element group 47: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_taken/$entry
      -- 
    convTransposeB_CP_4715_elements(47) <= convTransposeB_CP_4715_elements(52);
    -- CP-element group 48:  branch  place  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	215 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_body_done
      -- 
    convTransposeB_CP_4715_elements(48) <= convTransposeB_CP_4715_elements(215);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	61 
    -- CP-element group 49: 	82 
    -- CP-element group 49: 	103 
    -- CP-element group 49: 	124 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/back_edge_to_loop_body
      -- 
    convTransposeB_CP_4715_elements(49) <= convTransposeB_CP_4715_elements(46);
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	44 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	63 
    -- CP-element group 50: 	84 
    -- CP-element group 50: 	105 
    -- CP-element group 50: 	126 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/first_time_through_loop_body
      -- 
    convTransposeB_CP_4715_elements(50) <= convTransposeB_CP_4715_elements(44);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	57 
    -- CP-element group 51: 	58 
    -- CP-element group 51: 	76 
    -- CP-element group 51: 	77 
    -- CP-element group 51: 	97 
    -- CP-element group 51: 	98 
    -- CP-element group 51: 	118 
    -- CP-element group 51: 	119 
    -- CP-element group 51: 	156 
    -- CP-element group 51: 	157 
    -- CP-element group 51: 	167 
    -- CP-element group 51: 	169 
    -- CP-element group 51: 	186 
    -- CP-element group 51: 	214 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/$entry
      -- CP-element group 51: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/loop_body_start
      -- 
    -- Element group convTransposeB_CP_4715_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	213 
    -- CP-element group 52: 	214 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	47 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/condition_evaluated
      -- 
    condition_evaluated_5039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_5039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(52), ack => do_while_stmt_2007_branch_req_0); -- 
    convTransposeB_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(56) & convTransposeB_CP_4715_elements(213) & convTransposeB_CP_4715_elements(214);
      gj_convTransposeB_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	57 
    -- CP-element group 53: 	76 
    -- CP-element group 53: 	97 
    -- CP-element group 53: 	118 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53: 	99 
    -- CP-element group 53: 	120 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/aggregated_phi_sample_req
      -- CP-element group 53: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_sample_start__ps
      -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(57) & convTransposeB_CP_4715_elements(76) & convTransposeB_CP_4715_elements(97) & convTransposeB_CP_4715_elements(118) & convTransposeB_CP_4715_elements(56);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	59 
    -- CP-element group 54: 	79 
    -- CP-element group 54: 	100 
    -- CP-element group 54: 	121 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	183 
    -- CP-element group 54: 	187 
    -- CP-element group 54: 	191 
    -- CP-element group 54: 	195 
    -- CP-element group 54: 	199 
    -- CP-element group 54: 	203 
    -- CP-element group 54: 	207 
    -- CP-element group 54: 	215 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: 	76 
    -- CP-element group 54: 	97 
    -- CP-element group 54: 	118 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/aggregated_phi_sample_ack
      -- CP-element group 54: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_sample_completed_
      -- 
    convTransposeB_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(59) & convTransposeB_CP_4715_elements(79) & convTransposeB_CP_4715_elements(100) & convTransposeB_CP_4715_elements(121);
      gj_convTransposeB_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	77 
    -- CP-element group 55: 	98 
    -- CP-element group 55: 	119 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	80 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	122 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/aggregated_phi_update_req
      -- CP-element group 55: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_update_start__ps
      -- 
    convTransposeB_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(58) & convTransposeB_CP_4715_elements(77) & convTransposeB_CP_4715_elements(98) & convTransposeB_CP_4715_elements(119);
      gj_convTransposeB_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	81 
    -- CP-element group 56: 	102 
    -- CP-element group 56: 	123 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/aggregated_phi_update_ack
      -- 
    convTransposeB_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(60) & convTransposeB_CP_4715_elements(81) & convTransposeB_CP_4715_elements(102) & convTransposeB_CP_4715_elements(123);
      gj_convTransposeB_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	53 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_sample_start_
      -- 
    convTransposeB_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(54);
      gj_convTransposeB_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	153 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	55 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_update_start_
      -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(60) & convTransposeB_CP_4715_elements(153);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_sample_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: 	151 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_update_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	49 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_loopback_trigger
      -- 
    convTransposeB_CP_4715_elements(61) <= convTransposeB_CP_4715_elements(49);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_loopback_sample_req_ps
      -- 
    phi_stmt_2009_loopback_sample_req_5054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2009_loopback_sample_req_5054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(62), ack => phi_stmt_2009_req_0); -- 
    -- Element group convTransposeB_CP_4715_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	50 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_entry_trigger
      -- 
    convTransposeB_CP_4715_elements(63) <= convTransposeB_CP_4715_elements(50);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_entry_sample_req_ps
      -- 
    phi_stmt_2009_entry_sample_req_5057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2009_entry_sample_req_5057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(64), ack => phi_stmt_2009_req_1); -- 
    -- Element group convTransposeB_CP_4715_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2009_phi_mux_ack_ps
      -- 
    phi_stmt_2009_phi_mux_ack_5060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2009_ack_0, ack => convTransposeB_CP_4715_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_sample_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_update_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Sample/rr
      -- 
    rr_5073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(68), ack => type_cast_2012_inst_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(66) & convTransposeB_CP_4715_elements(70);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_update_start_
      -- CP-element group 69: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Update/cr
      -- 
    cr_5078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(69), ack => type_cast_2012_inst_req_1); -- 
    convTransposeB_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(67) & convTransposeB_CP_4715_elements(71);
      gj_convTransposeB_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Sample/ra
      -- 
    ra_5074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2012_inst_ack_0, ack => convTransposeB_CP_4715_elements(70)); -- 
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2012_Update/ca
      -- 
    ca_5079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2012_inst_ack_1, ack => convTransposeB_CP_4715_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_sample_completed_
      -- 
    -- Element group convTransposeB_CP_4715_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_update_start_
      -- 
    -- Element group convTransposeB_CP_4715_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_update_completed__ps
      -- 
    convTransposeB_CP_4715_elements(74) <= convTransposeB_CP_4715_elements(75);
    -- CP-element group 75:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_indvar_at_entry_2013_update_completed_
      -- 
    -- Element group convTransposeB_CP_4715_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeB_CP_4715_elements(73), ack => convTransposeB_CP_4715_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	51 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	54 
    -- CP-element group 76: 	185 
    -- CP-element group 76: 	189 
    -- CP-element group 76: 	193 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	53 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_sample_start_
      -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(185) & convTransposeB_CP_4715_elements(189) & convTransposeB_CP_4715_elements(193);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	51 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: 	141 
    -- CP-element group 77: 	184 
    -- CP-element group 77: 	192 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	55 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_update_start_
      -- 
    convTransposeB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(81) & convTransposeB_CP_4715_elements(141) & convTransposeB_CP_4715_elements(184) & convTransposeB_CP_4715_elements(192);
      gj_convTransposeB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	53 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_sample_start__ps
      -- 
    convTransposeB_CP_4715_elements(78) <= convTransposeB_CP_4715_elements(53);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	54 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_sample_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	55 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_update_start__ps
      -- 
    convTransposeB_CP_4715_elements(80) <= convTransposeB_CP_4715_elements(55);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	56 
    -- CP-element group 81: 	139 
    -- CP-element group 81: 	182 
    -- CP-element group 81: 	190 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_update_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	49 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_loopback_trigger
      -- 
    convTransposeB_CP_4715_elements(82) <= convTransposeB_CP_4715_elements(49);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_loopback_sample_req_ps
      -- 
    phi_stmt_2014_loopback_sample_req_5098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2014_loopback_sample_req_5098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(83), ack => phi_stmt_2014_req_1); -- 
    -- Element group convTransposeB_CP_4715_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	50 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_entry_trigger
      -- 
    convTransposeB_CP_4715_elements(84) <= convTransposeB_CP_4715_elements(50);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_entry_sample_req_ps
      -- 
    phi_stmt_2014_entry_sample_req_5101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2014_entry_sample_req_5101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(85), ack => phi_stmt_2014_req_0); -- 
    -- Element group convTransposeB_CP_4715_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_phi_mux_ack
      -- CP-element group 86: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2014_phi_mux_ack_ps
      -- 
    phi_stmt_2014_phi_mux_ack_5104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2014_ack_0, ack => convTransposeB_CP_4715_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_sample_start_
      -- 
    -- Element group convTransposeB_CP_4715_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_update_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_update_completed__ps
      -- 
    convTransposeB_CP_4715_elements(89) <= convTransposeB_CP_4715_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim2x_x1_at_entry_2016_update_completed_
      -- 
    -- Element group convTransposeB_CP_4715_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => convTransposeB_CP_4715_elements(88), ack => convTransposeB_CP_4715_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_sample_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_update_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_sample_start_
      -- 
    rr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(93), ack => type_cast_2018_inst_req_0); -- 
    convTransposeB_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(91) & convTransposeB_CP_4715_elements(95);
      gj_convTransposeB_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_update_start_
      -- 
    cr_5130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(94), ack => type_cast_2018_inst_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(92) & convTransposeB_CP_4715_elements(96);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_sample_completed__ps
      -- 
    ra_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_0, ack => convTransposeB_CP_4715_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2018_Update/ca
      -- 
    ca_5131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_1, ack => convTransposeB_CP_4715_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	51 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	54 
    -- CP-element group 97: 	197 
    -- CP-element group 97: 	201 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	53 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_sample_start_
      -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(197) & convTransposeB_CP_4715_elements(201);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	51 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: 	145 
    -- CP-element group 98: 	200 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	55 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_update_start_
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(102) & convTransposeB_CP_4715_elements(145) & convTransposeB_CP_4715_elements(200);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	53 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_sample_start__ps
      -- 
    convTransposeB_CP_4715_elements(99) <= convTransposeB_CP_4715_elements(53);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	54 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_sample_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_update_start__ps
      -- 
    convTransposeB_CP_4715_elements(101) <= convTransposeB_CP_4715_elements(55);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	56 
    -- CP-element group 102: 	143 
    -- CP-element group 102: 	198 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_update_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	49 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_loopback_trigger
      -- 
    convTransposeB_CP_4715_elements(103) <= convTransposeB_CP_4715_elements(49);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_loopback_sample_req
      -- 
    phi_stmt_2019_loopback_sample_req_5142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2019_loopback_sample_req_5142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(104), ack => phi_stmt_2019_req_1); -- 
    -- Element group convTransposeB_CP_4715_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	50 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_entry_trigger
      -- 
    convTransposeB_CP_4715_elements(105) <= convTransposeB_CP_4715_elements(50);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_entry_sample_req
      -- 
    phi_stmt_2019_entry_sample_req_5145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2019_entry_sample_req_5145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(106), ack => phi_stmt_2019_req_0); -- 
    -- Element group convTransposeB_CP_4715_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_phi_mux_ack_ps
      -- CP-element group 107: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2019_phi_mux_ack
      -- 
    phi_stmt_2019_phi_mux_ack_5148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2019_ack_0, ack => convTransposeB_CP_4715_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_sample_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_update_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_update_completed__ps
      -- 
    convTransposeB_CP_4715_elements(110) <= convTransposeB_CP_4715_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim1x_x1_at_entry_2021_update_completed_
      -- 
    -- Element group convTransposeB_CP_4715_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => convTransposeB_CP_4715_elements(109), ack => convTransposeB_CP_4715_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_sample_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_update_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_sample_start_
      -- 
    rr_5169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(114), ack => type_cast_2023_inst_req_0); -- 
    convTransposeB_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(112) & convTransposeB_CP_4715_elements(116);
      gj_convTransposeB_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_update_start_
      -- 
    cr_5174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(115), ack => type_cast_2023_inst_req_1); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(113) & convTransposeB_CP_4715_elements(117);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_sample_completed__ps
      -- 
    ra_5170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2023_inst_ack_0, ack => convTransposeB_CP_4715_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2023_update_completed__ps
      -- 
    ca_5175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2023_inst_ack_1, ack => convTransposeB_CP_4715_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	51 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	54 
    -- CP-element group 118: 	205 
    -- CP-element group 118: 	209 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	53 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_sample_start_
      -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(205) & convTransposeB_CP_4715_elements(209);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	51 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	149 
    -- CP-element group 119: 	208 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	55 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_update_start_
      -- 
    convTransposeB_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(123) & convTransposeB_CP_4715_elements(149) & convTransposeB_CP_4715_elements(208);
      gj_convTransposeB_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	53 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_sample_start__ps
      -- 
    convTransposeB_CP_4715_elements(120) <= convTransposeB_CP_4715_elements(53);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	54 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_sample_completed__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	55 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_update_start__ps
      -- 
    convTransposeB_CP_4715_elements(122) <= convTransposeB_CP_4715_elements(55);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	56 
    -- CP-element group 123: 	147 
    -- CP-element group 123: 	206 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	119 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_update_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_update_completed_
      -- 
    -- Element group convTransposeB_CP_4715_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	49 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_loopback_trigger
      -- 
    convTransposeB_CP_4715_elements(124) <= convTransposeB_CP_4715_elements(49);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_loopback_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_loopback_sample_req
      -- 
    phi_stmt_2024_loopback_sample_req_5186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2024_loopback_sample_req_5186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(125), ack => phi_stmt_2024_req_0); -- 
    -- Element group convTransposeB_CP_4715_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	50 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_entry_trigger
      -- 
    convTransposeB_CP_4715_elements(126) <= convTransposeB_CP_4715_elements(50);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_entry_sample_req_ps
      -- CP-element group 127: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_entry_sample_req
      -- 
    phi_stmt_2024_entry_sample_req_5189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2024_entry_sample_req_5189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(127), ack => phi_stmt_2024_req_1); -- 
    -- Element group convTransposeB_CP_4715_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_phi_mux_ack_ps
      -- CP-element group 128: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/phi_stmt_2024_phi_mux_ack
      -- 
    phi_stmt_2024_phi_mux_ack_5192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2024_ack_0, ack => convTransposeB_CP_4715_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_sample_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_update_start__ps
      -- 
    -- Element group convTransposeB_CP_4715_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_sample_start_
      -- 
    rr_5205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(131), ack => type_cast_2027_inst_req_0); -- 
    convTransposeB_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(129) & convTransposeB_CP_4715_elements(133);
      gj_convTransposeB_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_update_start_
      -- 
    cr_5210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(132), ack => type_cast_2027_inst_req_1); -- 
    convTransposeB_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(130) & convTransposeB_CP_4715_elements(134);
      gj_convTransposeB_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_sample_completed__ps
      -- 
    ra_5206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2027_inst_ack_0, ack => convTransposeB_CP_4715_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2027_update_completed__ps
      -- 
    ca_5211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2027_inst_ack_1, ack => convTransposeB_CP_4715_elements(134)); -- 
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Sample/req
      -- CP-element group 135: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_sample_start__ps
      -- 
    req_5223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(135), ack => input_dim0x_x1_at_entry_2002_2028_buf_req_0); -- 
    -- Element group convTransposeB_CP_4715_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Update/req
      -- CP-element group 136: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_update_start_
      -- CP-element group 136: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_update_start__ps
      -- 
    req_5228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(136), ack => input_dim0x_x1_at_entry_2002_2028_buf_req_1); -- 
    -- Element group convTransposeB_CP_4715_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_sample_completed__ps
      -- 
    ack_5224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_dim0x_x1_at_entry_2002_2028_buf_ack_0, ack => convTransposeB_CP_4715_elements(137)); -- 
    -- CP-element group 138:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Update/ack
      -- CP-element group 138: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/R_input_dim0x_x1_at_entry_2028_update_completed__ps
      -- 
    ack_5229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_dim0x_x1_at_entry_2002_2028_buf_ack_1, ack => convTransposeB_CP_4715_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	81 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_sample_start_
      -- 
    rr_5238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(139), ack => type_cast_2057_inst_req_0); -- 
    convTransposeB_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(81) & convTransposeB_CP_4715_elements(141);
      gj_convTransposeB_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: 	170 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_update_start_
      -- CP-element group 140: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Update/cr
      -- CP-element group 140: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Update/$entry
      -- 
    cr_5243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(140), ack => type_cast_2057_inst_req_1); -- 
    convTransposeB_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(142) & convTransposeB_CP_4715_elements(170);
      gj_convTransposeB_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	77 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Sample/ra
      -- 
    ra_5239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2057_inst_ack_0, ack => convTransposeB_CP_4715_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	168 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2057_Update/ca
      -- 
    ca_5244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2057_inst_ack_1, ack => convTransposeB_CP_4715_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	102 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_sample_start_
      -- 
    rr_5252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(143), ack => type_cast_2061_inst_req_0); -- 
    convTransposeB_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(102) & convTransposeB_CP_4715_elements(145);
      gj_convTransposeB_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: 	170 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_update_start_
      -- 
    cr_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(144), ack => type_cast_2061_inst_req_1); -- 
    convTransposeB_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(146) & convTransposeB_CP_4715_elements(170);
      gj_convTransposeB_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	98 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_sample_completed_
      -- 
    ra_5253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_0, ack => convTransposeB_CP_4715_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	168 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2061_update_completed_
      -- 
    ca_5258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_1, ack => convTransposeB_CP_4715_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	123 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_sample_start_
      -- 
    rr_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(147), ack => type_cast_2065_inst_req_0); -- 
    convTransposeB_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(123) & convTransposeB_CP_4715_elements(149);
      gj_convTransposeB_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: 	170 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Update/cr
      -- CP-element group 148: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_update_start_
      -- 
    cr_5271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(148), ack => type_cast_2065_inst_req_1); -- 
    convTransposeB_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(150) & convTransposeB_CP_4715_elements(170);
      gj_convTransposeB_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	119 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_sample_completed_
      -- 
    ra_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_0, ack => convTransposeB_CP_4715_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	168 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2065_update_completed_
      -- 
    ca_5272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2065_inst_ack_1, ack => convTransposeB_CP_4715_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	60 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_sample_start_
      -- 
    rr_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(151), ack => type_cast_2089_inst_req_0); -- 
    convTransposeB_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(60) & convTransposeB_CP_4715_elements(153);
      gj_convTransposeB_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: 	158 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Update/cr
      -- CP-element group 152: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_update_start_
      -- CP-element group 152: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Update/$entry
      -- 
    cr_5285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(152), ack => type_cast_2089_inst_req_1); -- 
    convTransposeB_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(154) & convTransposeB_CP_4715_elements(158);
      gj_convTransposeB_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	58 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_sample_completed_
      -- 
    ra_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2089_inst_ack_0, ack => convTransposeB_CP_4715_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	158 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (16) 
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_resized_1
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2089_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_scaled_1
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_scale_1/scale_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_scale_1/scale_rename_req
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_scale_1/$exit
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_scale_1/$entry
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_resize_1/index_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_resize_1/index_resize_req
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_resize_1/$exit
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_resize_1/$entry
      -- CP-element group 154: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_index_computed_1
      -- 
    ca_5286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2089_inst_ack_1, ack => convTransposeB_CP_4715_elements(154)); -- 
    req_5311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(154), ack => array_obj_ref_2095_index_offset_req_0); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	160 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	160 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_request/req
      -- CP-element group 155: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_request/$entry
      -- 
    req_5326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(155), ack => addr_of_2096_final_reg_req_0); -- 
    convTransposeB_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(159) & convTransposeB_CP_4715_elements(160);
      gj_convTransposeB_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	51 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	164 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_update_start_
      -- CP-element group 156: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_complete/req
      -- 
    req_5331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(156), ack => addr_of_2096_final_reg_req_1); -- 
    convTransposeB_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(161) & convTransposeB_CP_4715_elements(164);
      gj_convTransposeB_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	51 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Update/req
      -- CP-element group 157: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_update_start
      -- 
    req_5316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(157), ack => array_obj_ref_2095_index_offset_req_1); -- 
    convTransposeB_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(159) & convTransposeB_CP_4715_elements(160);
      gj_convTransposeB_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	215 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	152 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Sample/ack
      -- CP-element group 158: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_sample_complete
      -- 
    ack_5312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2095_index_offset_ack_0, ack => convTransposeB_CP_4715_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (8) 
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_offset_calculated
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_base_plus_offset/sum_rename_req
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_base_plus_offset/sum_rename_ack
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_base_plus_offset/$entry
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_base_plus_offset/$exit
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_root_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Update/ack
      -- CP-element group 159: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2095_final_index_sum_regn_Update/$exit
      -- 
    ack_5317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2095_index_offset_ack_1, ack => convTransposeB_CP_4715_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_request/ack
      -- CP-element group 160: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_request/$exit
      -- 
    ack_5327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2096_final_reg_ack_0, ack => convTransposeB_CP_4715_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (19) 
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_addr_resize/base_resize_ack
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_addr_resize/base_resize_req
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_complete/ack
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_complete/$exit
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_word_addrgen/root_register_req
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_address_resized
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2096_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_word_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_root_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_addr_resize/$exit
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_addr_resize/$entry
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_word_addrgen/root_register_ack
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_word_addrgen/$exit
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_word_addrgen/$entry
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_plus_offset/sum_rename_ack
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_plus_offset/sum_rename_req
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_plus_offset/$exit
      -- CP-element group 161: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_base_plus_offset/$entry
      -- 
    ack_5332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2096_final_reg_ack_1, ack => convTransposeB_CP_4715_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/word_access_start/word_0/rr
      -- CP-element group 162: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/word_access_start/$entry
      -- 
    rr_5365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(162), ack => ptr_deref_2100_load_0_req_0); -- 
    convTransposeB_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(161) & convTransposeB_CP_4715_elements(164);
      gj_convTransposeB_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: 	180 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_update_start_
      -- 
    cr_5376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(163), ack => ptr_deref_2100_load_0_req_1); -- 
    convTransposeB_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(165) & convTransposeB_CP_4715_elements(180);
      gj_convTransposeB_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/word_access_start/word_0/ra
      -- CP-element group 164: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/word_access_start/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Sample/word_access_start/$exit
      -- 
    ra_5366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2100_load_0_ack_0, ack => convTransposeB_CP_4715_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	178 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (9) 
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/ptr_deref_2100_Merge/$entry
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/word_access_complete/word_0/ca
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/word_access_complete/word_0/$exit
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/ptr_deref_2100_Merge/$exit
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/ptr_deref_2100_Merge/merge_req
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/word_access_complete/$exit
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2100_Update/ptr_deref_2100_Merge/merge_ack
      -- 
    ca_5377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2100_load_0_ack_1, ack => convTransposeB_CP_4715_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	171 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	172 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	172 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_request/req
      -- CP-element group 166: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_request/$entry
      -- CP-element group 166: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_sample_start_
      -- 
    req_5422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(166), ack => addr_of_2119_final_reg_req_0); -- 
    convTransposeB_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(171) & convTransposeB_CP_4715_elements(172);
      gj_convTransposeB_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	51 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	173 
    -- CP-element group 167: 	176 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	173 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_complete/req
      -- CP-element group 167: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_update_start_
      -- 
    req_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(167), ack => addr_of_2119_final_reg_req_1); -- 
    convTransposeB_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(173) & convTransposeB_CP_4715_elements(176);
      gj_convTransposeB_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	142 
    -- CP-element group 168: 	146 
    -- CP-element group 168: 	150 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (13) 
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Sample/req
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_scale_1/scale_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_scale_1/scale_rename_req
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_scale_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_scale_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_resize_1/index_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_resize_1/index_resize_req
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_resize_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_resize_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_computed_1
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_scaled_1
      -- CP-element group 168: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_index_resized_1
      -- 
    req_5407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(168), ack => array_obj_ref_2118_index_offset_req_0); -- 
    convTransposeB_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(142) & convTransposeB_CP_4715_elements(146) & convTransposeB_CP_4715_elements(150);
      gj_convTransposeB_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	51 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Update/req
      -- CP-element group 169: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_update_start
      -- 
    req_5412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(169), ack => array_obj_ref_2118_index_offset_req_1); -- 
    convTransposeB_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(171) & convTransposeB_CP_4715_elements(172);
      gj_convTransposeB_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	215 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	140 
    -- CP-element group 170: 	144 
    -- CP-element group 170: 	148 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Sample/ack
      -- CP-element group 170: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_sample_complete
      -- 
    ack_5408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2118_index_offset_ack_0, ack => convTransposeB_CP_4715_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	166 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (8) 
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_base_plus_offset/sum_rename_ack
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/array_obj_ref_2118_root_address_calculated
      -- 
    ack_5413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2118_index_offset_ack_1, ack => convTransposeB_CP_4715_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_request/ack
      -- CP-element group 172: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_request/$exit
      -- CP-element group 172: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_sample_completed_
      -- 
    ack_5423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2119_final_reg_ack_0, ack => convTransposeB_CP_4715_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	167 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	167 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_complete/ack
      -- CP-element group 173: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/addr_of_2119_update_completed_
      -- 
    ack_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2119_final_reg_ack_1, ack => convTransposeB_CP_4715_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Sample/req
      -- CP-element group 174: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_sample_start_
      -- 
    req_5436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(174), ack => W_arrayidx86_2106_delayed_6_0_2121_inst_req_0); -- 
    convTransposeB_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(173) & convTransposeB_CP_4715_elements(176);
      gj_convTransposeB_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: 	180 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Update/req
      -- 
    req_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(175), ack => W_arrayidx86_2106_delayed_6_0_2121_inst_req_1); -- 
    convTransposeB_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(177) & convTransposeB_CP_4715_elements(180);
      gj_convTransposeB_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	167 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Sample/ack
      -- 
    ack_5437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx86_2106_delayed_6_0_2121_inst_ack_0, ack => convTransposeB_CP_4715_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (19) 
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_address_resized
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_addr_resize/$entry
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_addr_resize/base_resize_req
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_addr_resize/$exit
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_word_addrgen/root_register_ack
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_word_addrgen/root_register_req
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_word_addrgen/$exit
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_word_addrgen/$entry
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_root_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_plus_offset/sum_rename_ack
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_plus_offset/sum_rename_req
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_plus_offset/$exit
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_plus_offset/$entry
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_word_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Update/ack
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2123_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_base_addr_resize/base_resize_ack
      -- 
    ack_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx86_2106_delayed_6_0_2121_inst_ack_1, ack => convTransposeB_CP_4715_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	165 
    -- CP-element group 178: 	177 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/word_access_start/word_0/$entry
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/word_access_start/word_0/rr
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/ptr_deref_2125_Split/$exit
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/ptr_deref_2125_Split/split_ack
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/ptr_deref_2125_Split/$entry
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/ptr_deref_2125_Split/split_req
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/word_access_start/$entry
      -- 
    rr_5480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(178), ack => ptr_deref_2125_store_0_req_0); -- 
    convTransposeB_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(165) & convTransposeB_CP_4715_elements(177) & convTransposeB_CP_4715_elements(180);
      gj_convTransposeB_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (5) 
      -- CP-element group 179: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/word_access_complete/word_0/cr
      -- CP-element group 179: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/word_access_complete/word_0/$entry
      -- CP-element group 179: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/word_access_complete/$entry
      -- CP-element group 179: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_update_start_
      -- 
    cr_5491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(179), ack => ptr_deref_2125_store_0_req_1); -- 
    convTransposeB_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeB_CP_4715_elements(181);
      gj_convTransposeB_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	163 
    -- CP-element group 180: 	175 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/word_access_start/word_0/$exit
      -- CP-element group 180: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/word_access_start/word_0/ra
      -- CP-element group 180: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Sample/word_access_start/$exit
      -- CP-element group 180: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_sample_completed_
      -- 
    ra_5481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2125_store_0_ack_0, ack => convTransposeB_CP_4715_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	215 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/word_access_complete/word_0/ca
      -- CP-element group 181: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/word_access_complete/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_Update/word_access_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/ptr_deref_2125_update_completed_
      -- 
    ca_5492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2125_store_0_ack_1, ack => convTransposeB_CP_4715_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	81 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Sample/rr
      -- 
    rr_5500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(182), ack => type_cast_2130_inst_req_0); -- 
    convTransposeB_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(81) & convTransposeB_CP_4715_elements(184);
      gj_convTransposeB_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	54 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: 	196 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Update/$entry
      -- 
    cr_5505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(183), ack => type_cast_2130_inst_req_1); -- 
    convTransposeB_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(185) & convTransposeB_CP_4715_elements(196);
      gj_convTransposeB_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	77 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Sample/ra
      -- 
    ra_5501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2130_inst_ack_0, ack => convTransposeB_CP_4715_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	194 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	76 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2130_update_completed_
      -- 
    ca_5506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2130_inst_ack_1, ack => convTransposeB_CP_4715_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	51 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Sample/rr
      -- 
    rr_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(186), ack => type_cast_2134_inst_req_0); -- 
    convTransposeB_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(51) & convTransposeB_CP_4715_elements(188);
      gj_convTransposeB_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	54 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	189 
    -- CP-element group 187: 	196 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Update/cr
      -- 
    cr_5519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(187), ack => type_cast_2134_inst_req_1); -- 
    convTransposeB_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(189) & convTransposeB_CP_4715_elements(196);
      gj_convTransposeB_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Sample/ra
      -- 
    ra_5515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2134_inst_ack_0, ack => convTransposeB_CP_4715_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	194 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	76 
    -- CP-element group 189: 	187 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2134_Update/ca
      -- 
    ca_5520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2134_inst_ack_1, ack => convTransposeB_CP_4715_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	81 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Sample/req
      -- 
    req_5528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(190), ack => W_add101_2129_delayed_1_0_2148_inst_req_0); -- 
    convTransposeB_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(81) & convTransposeB_CP_4715_elements(192);
      gj_convTransposeB_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	54 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_update_start_
      -- CP-element group 191: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Update/req
      -- 
    req_5533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(191), ack => W_add101_2129_delayed_1_0_2148_inst_req_1); -- 
    convTransposeB_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(193);
      gj_convTransposeB_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	77 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Sample/ack
      -- 
    ack_5529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add101_2129_delayed_1_0_2148_inst_ack_0, ack => convTransposeB_CP_4715_elements(192)); -- 
    -- CP-element group 193:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	215 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	76 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2150_Update/ack
      -- 
    ack_5534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add101_2129_delayed_1_0_2148_inst_ack_1, ack => convTransposeB_CP_4715_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	185 
    -- CP-element group 194: 	189 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Sample/rr
      -- 
    rr_5542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(194), ack => type_cast_2160_inst_req_0); -- 
    convTransposeB_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(185) & convTransposeB_CP_4715_elements(189) & convTransposeB_CP_4715_elements(196);
      gj_convTransposeB_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	54 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: 	204 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Update/cr
      -- 
    cr_5547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(195), ack => type_cast_2160_inst_req_1); -- 
    convTransposeB_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(197) & convTransposeB_CP_4715_elements(204);
      gj_convTransposeB_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	183 
    -- CP-element group 196: 	187 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Sample/ra
      -- 
    ra_5543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2160_inst_ack_0, ack => convTransposeB_CP_4715_elements(196)); -- 
    -- CP-element group 197:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	202 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	97 
    -- CP-element group 197: 	195 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2160_Update/ca
      -- 
    ca_5548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2160_inst_ack_1, ack => convTransposeB_CP_4715_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	102 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Sample/req
      -- 
    req_5556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(198), ack => W_input_dim1x_x1_2146_delayed_2_0_2168_inst_req_0); -- 
    convTransposeB_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(102) & convTransposeB_CP_4715_elements(200);
      gj_convTransposeB_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	54 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	201 
    -- CP-element group 199: 	204 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_update_start_
      -- CP-element group 199: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Update/req
      -- 
    req_5561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(199), ack => W_input_dim1x_x1_2146_delayed_2_0_2168_inst_req_1); -- 
    convTransposeB_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(201) & convTransposeB_CP_4715_elements(204);
      gj_convTransposeB_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	98 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Sample/ack
      -- 
    ack_5557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_2146_delayed_2_0_2168_inst_ack_0, ack => convTransposeB_CP_4715_elements(200)); -- 
    -- CP-element group 201:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	97 
    -- CP-element group 201: 	199 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2170_Update/ack
      -- 
    ack_5562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_2146_delayed_2_0_2168_inst_ack_1, ack => convTransposeB_CP_4715_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	197 
    -- CP-element group 202: 	201 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Sample/rr
      -- 
    rr_5570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(202), ack => type_cast_2183_inst_req_0); -- 
    convTransposeB_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(197) & convTransposeB_CP_4715_elements(201) & convTransposeB_CP_4715_elements(204);
      gj_convTransposeB_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	54 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: 	212 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_update_start_
      -- CP-element group 203: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Update/cr
      -- 
    cr_5575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(203), ack => type_cast_2183_inst_req_1); -- 
    convTransposeB_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(205) & convTransposeB_CP_4715_elements(212);
      gj_convTransposeB_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	195 
    -- CP-element group 204: 	199 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Sample/ra
      -- 
    ra_5571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2183_inst_ack_0, ack => convTransposeB_CP_4715_elements(204)); -- 
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	210 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	118 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2183_Update/ca
      -- 
    ca_5576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2183_inst_ack_1, ack => convTransposeB_CP_4715_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	123 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Sample/req
      -- 
    req_5584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(206), ack => W_input_dim0x_x1_2160_delayed_3_0_2185_inst_req_0); -- 
    convTransposeB_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(123) & convTransposeB_CP_4715_elements(208);
      gj_convTransposeB_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	54 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: 	212 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_update_start_
      -- CP-element group 207: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Update/req
      -- 
    req_5589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(207), ack => W_input_dim0x_x1_2160_delayed_3_0_2185_inst_req_1); -- 
    convTransposeB_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(209) & convTransposeB_CP_4715_elements(212);
      gj_convTransposeB_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	119 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Sample/ack
      -- 
    ack_5585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_2160_delayed_3_0_2185_inst_ack_0, ack => convTransposeB_CP_4715_elements(208)); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	118 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/assign_stmt_2187_Update/ack
      -- 
    ack_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_2160_delayed_3_0_2185_inst_ack_1, ack => convTransposeB_CP_4715_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	205 
    -- CP-element group 210: 	209 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Sample/rr
      -- 
    rr_5598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(210), ack => type_cast_2202_inst_req_0); -- 
    convTransposeB_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(205) & convTransposeB_CP_4715_elements(209) & convTransposeB_CP_4715_elements(212);
      gj_convTransposeB_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_update_start_
      -- CP-element group 211: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Update/cr
      -- 
    cr_5603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(211), ack => type_cast_2202_inst_req_1); -- 
    convTransposeB_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeB_CP_4715_elements(213);
      gj_convTransposeB_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	203 
    -- CP-element group 212: 	207 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Sample/ra
      -- 
    ra_5599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2202_inst_ack_0, ack => convTransposeB_CP_4715_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	52 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/type_cast_2202_Update/ca
      -- 
    ca_5604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2202_inst_ack_1, ack => convTransposeB_CP_4715_elements(213)); -- 
    -- CP-element group 214:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	51 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	52 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convTransposeB_CP_4715_elements(214) is a control-delay.
    cp_element_214_delay: control_delay_element  generic map(name => " 214_delay", delay_value => 1)  port map(req => convTransposeB_CP_4715_elements(51), ack => convTransposeB_CP_4715_elements(214), clk => clk, reset =>reset);
    -- CP-element group 215:  join  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	54 
    -- CP-element group 215: 	158 
    -- CP-element group 215: 	170 
    -- CP-element group 215: 	181 
    -- CP-element group 215: 	193 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	48 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_1865/do_while_stmt_2007/do_while_stmt_2007_loop_body/$exit
      -- 
    convTransposeB_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(54) & convTransposeB_CP_4715_elements(158) & convTransposeB_CP_4715_elements(170) & convTransposeB_CP_4715_elements(181) & convTransposeB_CP_4715_elements(193);
      gj_convTransposeB_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_exit/$exit
      -- CP-element group 216: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_exit/ack
      -- 
    ack_5609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2007_branch_ack_0, ack => convTransposeB_CP_4715_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	47 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_taken/$exit
      -- CP-element group 217: 	 branch_block_stmt_1865/do_while_stmt_2007/loop_taken/ack
      -- 
    ack_5613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2007_branch_ack_1, ack => convTransposeB_CP_4715_elements(217)); -- 
    -- CP-element group 218:  transition  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	1 
    -- CP-element group 218:  members (1) 
      -- CP-element group 218: 	 branch_block_stmt_1865/do_while_stmt_2007/$exit
      -- 
    convTransposeB_CP_4715_elements(218) <= convTransposeB_CP_4715_elements(45);
    -- CP-element group 219:  merge  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	1 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (15) 
      -- CP-element group 219: 	 branch_block_stmt_1865/assign_stmt_2230__entry__
      -- CP-element group 219: 	 branch_block_stmt_1865/merge_stmt_2225__exit__
      -- CP-element group 219: 	 branch_block_stmt_1865/if_stmt_2221_if_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_1865/if_stmt_2221_if_link/if_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_1865/whilex_xbody_whilex_xend
      -- CP-element group 219: 	 branch_block_stmt_1865/assign_stmt_2230/$entry
      -- CP-element group 219: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Sample/req
      -- CP-element group 219: 	 branch_block_stmt_1865/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_1865/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_1865/merge_stmt_2225_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_1865/merge_stmt_2225_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_1865/merge_stmt_2225_PhiAck/$exit
      -- CP-element group 219: 	 branch_block_stmt_1865/merge_stmt_2225_PhiAck/dummy
      -- 
    if_choice_transition_5627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2221_branch_ack_1, ack => convTransposeB_CP_4715_elements(219)); -- 
    req_5643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(219), ack => WPIPE_Block1_done_2227_inst_req_0); -- 
    -- CP-element group 220:  merge  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	1 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_1865/merge_stmt_2225__entry__
      -- CP-element group 220: 	 branch_block_stmt_1865/if_stmt_2221__exit__
      -- CP-element group 220: 	 branch_block_stmt_1865/if_stmt_2221_else_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_1865/if_stmt_2221_else_link/else_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_1865/merge_stmt_2225_dead_link/$entry
      -- 
    else_choice_transition_5631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2221_branch_ack_0, ack => convTransposeB_CP_4715_elements(220)); -- 
    -- CP-element group 221:  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_update_start_
      -- CP-element group 221: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Sample/ack
      -- CP-element group 221: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Update/req
      -- 
    ack_5644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2227_inst_ack_0, ack => convTransposeB_CP_4715_elements(221)); -- 
    req_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(221), ack => WPIPE_Block1_done_2227_inst_req_1); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (16) 
      -- CP-element group 222: 	 branch_block_stmt_1865/merge_stmt_2232__exit__
      -- CP-element group 222: 	 branch_block_stmt_1865/return__
      -- CP-element group 222: 	 branch_block_stmt_1865/assign_stmt_2230__exit__
      -- CP-element group 222: 	 $exit
      -- CP-element group 222: 	 branch_block_stmt_1865/branch_block_stmt_1865__exit__
      -- CP-element group 222: 	 branch_block_stmt_1865/$exit
      -- CP-element group 222: 	 branch_block_stmt_1865/assign_stmt_2230/$exit
      -- CP-element group 222: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_1865/assign_stmt_2230/WPIPE_Block1_done_2227_Update/ack
      -- CP-element group 222: 	 branch_block_stmt_1865/return___PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_1865/return___PhiReq/$exit
      -- CP-element group 222: 	 branch_block_stmt_1865/merge_stmt_2232_PhiReqMerge
      -- CP-element group 222: 	 branch_block_stmt_1865/merge_stmt_2232_PhiAck/$entry
      -- CP-element group 222: 	 branch_block_stmt_1865/merge_stmt_2232_PhiAck/$exit
      -- CP-element group 222: 	 branch_block_stmt_1865/merge_stmt_2232_PhiAck/dummy
      -- 
    ack_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2227_inst_ack_1, ack => convTransposeB_CP_4715_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	43 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Sample/ra
      -- 
    ra_5669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2005_inst_ack_0, ack => convTransposeB_CP_4715_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	43 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/Update/ca
      -- 
    ca_5674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2005_inst_ack_1, ack => convTransposeB_CP_4715_elements(224)); -- 
    -- CP-element group 225:  join  transition  place  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (8) 
      -- CP-element group 225: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/$exit
      -- CP-element group 225: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/$exit
      -- CP-element group 225: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/$exit
      -- CP-element group 225: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/$exit
      -- CP-element group 225: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_sources/type_cast_2005/SplitProtocol/$exit
      -- CP-element group 225: 	 branch_block_stmt_1865/entry_whilex_xbody_PhiReq/phi_stmt_2002/phi_stmt_2002_req
      -- CP-element group 225: 	 branch_block_stmt_1865/merge_stmt_1986_PhiReqMerge
      -- CP-element group 225: 	 branch_block_stmt_1865/merge_stmt_1986_PhiAck/$entry
      -- 
    phi_stmt_2002_req_5675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2002_req_5675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4715_elements(225), ack => phi_stmt_2002_req_0); -- 
    convTransposeB_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4715_elements(223) & convTransposeB_CP_4715_elements(224);
      gj_convTransposeB_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4715_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  transition  place  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	44 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_1865/do_while_stmt_2007__entry__
      -- CP-element group 226: 	 branch_block_stmt_1865/merge_stmt_1986__exit__
      -- CP-element group 226: 	 branch_block_stmt_1865/merge_stmt_1986_PhiAck/$exit
      -- CP-element group 226: 	 branch_block_stmt_1865/merge_stmt_1986_PhiAck/phi_stmt_2002_ack
      -- 
    phi_stmt_2002_ack_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2002_ack_0, ack => convTransposeB_CP_4715_elements(226)); -- 
    convTransposeB_do_while_stmt_2007_terminator_5614: loop_terminator -- 
      generic map (name => " convTransposeB_do_while_stmt_2007_terminator_5614", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convTransposeB_CP_4715_elements(48),loop_continue => convTransposeB_CP_4715_elements(217),loop_terminate => convTransposeB_CP_4715_elements(216),loop_back => convTransposeB_CP_4715_elements(46),loop_exit => convTransposeB_CP_4715_elements(45),clk => clk, reset => reset); -- 
    phi_stmt_2009_phi_seq_5088_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeB_CP_4715_elements(61);
      convTransposeB_CP_4715_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeB_CP_4715_elements(70);
      convTransposeB_CP_4715_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeB_CP_4715_elements(71);
      convTransposeB_CP_4715_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeB_CP_4715_elements(63);
      convTransposeB_CP_4715_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeB_CP_4715_elements(72);
      convTransposeB_CP_4715_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeB_CP_4715_elements(74);
      convTransposeB_CP_4715_elements(64) <= phi_mux_reqs(1);
      phi_stmt_2009_phi_seq_5088 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2009_phi_seq_5088") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeB_CP_4715_elements(53), 
          phi_sample_ack => convTransposeB_CP_4715_elements(59), 
          phi_update_req => convTransposeB_CP_4715_elements(55), 
          phi_update_ack => convTransposeB_CP_4715_elements(60), 
          phi_mux_ack => convTransposeB_CP_4715_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2014_phi_seq_5132_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeB_CP_4715_elements(84);
      convTransposeB_CP_4715_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeB_CP_4715_elements(87);
      convTransposeB_CP_4715_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeB_CP_4715_elements(89);
      convTransposeB_CP_4715_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeB_CP_4715_elements(82);
      convTransposeB_CP_4715_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeB_CP_4715_elements(95);
      convTransposeB_CP_4715_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeB_CP_4715_elements(96);
      convTransposeB_CP_4715_elements(83) <= phi_mux_reqs(1);
      phi_stmt_2014_phi_seq_5132 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2014_phi_seq_5132") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeB_CP_4715_elements(78), 
          phi_sample_ack => convTransposeB_CP_4715_elements(79), 
          phi_update_req => convTransposeB_CP_4715_elements(80), 
          phi_update_ack => convTransposeB_CP_4715_elements(81), 
          phi_mux_ack => convTransposeB_CP_4715_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2019_phi_seq_5176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeB_CP_4715_elements(105);
      convTransposeB_CP_4715_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeB_CP_4715_elements(108);
      convTransposeB_CP_4715_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeB_CP_4715_elements(110);
      convTransposeB_CP_4715_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeB_CP_4715_elements(103);
      convTransposeB_CP_4715_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeB_CP_4715_elements(116);
      convTransposeB_CP_4715_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeB_CP_4715_elements(117);
      convTransposeB_CP_4715_elements(104) <= phi_mux_reqs(1);
      phi_stmt_2019_phi_seq_5176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2019_phi_seq_5176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeB_CP_4715_elements(99), 
          phi_sample_ack => convTransposeB_CP_4715_elements(100), 
          phi_update_req => convTransposeB_CP_4715_elements(101), 
          phi_update_ack => convTransposeB_CP_4715_elements(102), 
          phi_mux_ack => convTransposeB_CP_4715_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2024_phi_seq_5230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeB_CP_4715_elements(124);
      convTransposeB_CP_4715_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeB_CP_4715_elements(133);
      convTransposeB_CP_4715_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeB_CP_4715_elements(134);
      convTransposeB_CP_4715_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeB_CP_4715_elements(126);
      convTransposeB_CP_4715_elements(135)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeB_CP_4715_elements(137);
      convTransposeB_CP_4715_elements(136)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeB_CP_4715_elements(138);
      convTransposeB_CP_4715_elements(127) <= phi_mux_reqs(1);
      phi_stmt_2024_phi_seq_5230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2024_phi_seq_5230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeB_CP_4715_elements(120), 
          phi_sample_ack => convTransposeB_CP_4715_elements(121), 
          phi_update_req => convTransposeB_CP_4715_elements(122), 
          phi_update_ack => convTransposeB_CP_4715_elements(123), 
          phi_mux_ack => convTransposeB_CP_4715_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_5040_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convTransposeB_CP_4715_elements(49);
        preds(1)  <= convTransposeB_CP_4715_elements(50);
        entry_tmerge_5040 : transition_merge -- 
          generic map(name => " entry_tmerge_5040")
          port map (preds => preds, symbol_out => convTransposeB_CP_4715_elements(51));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_2220_wire : std_logic_vector(0 downto 0);
    signal R_idxprom85_2117_resized : std_logic_vector(13 downto 0);
    signal R_idxprom85_2117_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2094_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2094_scaled : std_logic_vector(13 downto 0);
    signal add101_2129_delayed_1_0_2150 : std_logic_vector(15 downto 0);
    signal add101_2147 : std_logic_vector(15 downto 0);
    signal add45_1939 : std_logic_vector(15 downto 0);
    signal add58_1950 : std_logic_vector(15 downto 0);
    signal add77_2076 : std_logic_vector(63 downto 0);
    signal add79_2086 : std_logic_vector(63 downto 0);
    signal add_1917 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2034 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2095_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2095_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2118_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2118_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2118_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2118_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2118_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2118_root_address : std_logic_vector(13 downto 0);
    signal arrayidx81_2097 : std_logic_vector(31 downto 0);
    signal arrayidx86_2106_delayed_6_0_2123 : std_logic_vector(31 downto 0);
    signal arrayidx86_2120 : std_logic_vector(31 downto 0);
    signal call11_1886 : std_logic_vector(15 downto 0);
    signal call13_1889 : std_logic_vector(15 downto 0);
    signal call14_1892 : std_logic_vector(15 downto 0);
    signal call15_1895 : std_logic_vector(15 downto 0);
    signal call16_1908 : std_logic_vector(15 downto 0);
    signal call18_1920 : std_logic_vector(15 downto 0);
    signal call1_1871 : std_logic_vector(15 downto 0);
    signal call20_1923 : std_logic_vector(15 downto 0);
    signal call22_1926 : std_logic_vector(15 downto 0);
    signal call3_1874 : std_logic_vector(15 downto 0);
    signal call5_1877 : std_logic_vector(15 downto 0);
    signal call7_1880 : std_logic_vector(15 downto 0);
    signal call9_1883 : std_logic_vector(15 downto 0);
    signal call_1868 : std_logic_vector(15 downto 0);
    signal cmp109_2180 : std_logic_vector(0 downto 0);
    signal cmp121_2208 : std_logic_vector(0 downto 0);
    signal cmp_2141 : std_logic_vector(0 downto 0);
    signal conv116_2203 : std_logic_vector(31 downto 0);
    signal conv119_1978 : std_logic_vector(31 downto 0);
    signal conv17_1912 : std_logic_vector(31 downto 0);
    signal conv65_2058 : std_logic_vector(63 downto 0);
    signal conv68_1959 : std_logic_vector(63 downto 0);
    signal conv70_2062 : std_logic_vector(63 downto 0);
    signal conv73_1963 : std_logic_vector(63 downto 0);
    signal conv75_2066 : std_logic_vector(63 downto 0);
    signal conv95_2131 : std_logic_vector(31 downto 0);
    signal conv97_1974 : std_logic_vector(31 downto 0);
    signal conv_1899 : std_logic_vector(31 downto 0);
    signal iNsTr_18_2161 : std_logic_vector(15 downto 0);
    signal idxprom85_2113 : std_logic_vector(63 downto 0);
    signal idxprom_2090 : std_logic_vector(63 downto 0);
    signal inc113_2184 : std_logic_vector(15 downto 0);
    signal inc113x_xinput_dim0x_x1_2192 : std_logic_vector(15 downto 0);
    signal inc_2167 : std_logic_vector(15 downto 0);
    signal indvar_2009 : std_logic_vector(31 downto 0);
    signal indvar_at_entry_1987 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2214 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1_2024 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_2160_delayed_3_0_2187 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_2002 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_2002_2028_buffered : std_logic_vector(15 downto 0);
    signal input_dim1x_x0_2175 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2019 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2146_delayed_2_0_2170 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_at_entry_1997 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2199 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0_2157 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2014 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_at_entry_1992 : std_logic_vector(15 downto 0);
    signal mul54_2049 : std_logic_vector(15 downto 0);
    signal mul76_2071 : std_logic_vector(63 downto 0);
    signal mul78_2081 : std_logic_vector(63 downto 0);
    signal mul_2039 : std_logic_vector(15 downto 0);
    signal ptr_deref_2100_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2100_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2125_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2125_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2125_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2125_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2125_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2125_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1905 : std_logic_vector(31 downto 0);
    signal shr120135_1984 : std_logic_vector(31 downto 0);
    signal shr134_1933 : std_logic_vector(15 downto 0);
    signal shr84_2107 : std_logic_vector(63 downto 0);
    signal sub48_2044 : std_logic_vector(15 downto 0);
    signal sub61_1955 : std_logic_vector(15 downto 0);
    signal sub62_2054 : std_logic_vector(15 downto 0);
    signal sub91_1969 : std_logic_vector(15 downto 0);
    signal sub_1944 : std_logic_vector(15 downto 0);
    signal tmp82_2101 : std_logic_vector(63 downto 0);
    signal type_cast_1903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1931_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1937_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1948_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1967_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1972_wire : std_logic_vector(31 downto 0);
    signal type_cast_1982_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2005_wire : std_logic_vector(15 downto 0);
    signal type_cast_2012_wire : std_logic_vector(31 downto 0);
    signal type_cast_2018_wire : std_logic_vector(15 downto 0);
    signal type_cast_2023_wire : std_logic_vector(15 downto 0);
    signal type_cast_2027_wire : std_logic_vector(15 downto 0);
    signal type_cast_2105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2111_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2118_2118_delayed_2_0_2135 : std_logic_vector(31 downto 0);
    signal type_cast_2138_wire : std_logic_vector(31 downto 0);
    signal type_cast_2145_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2155_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2165_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2196_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2212_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2229_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_whilex_xend_taken_2217 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_2095_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2095_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2095_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2095_resized_base_address <= "00000000000000";
    array_obj_ref_2118_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2118_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2118_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2118_resized_base_address <= "00000000000000";
    indvar_at_entry_1987 <= "00000000000000000000000000000000";
    input_dim1x_x1_at_entry_1997 <= "0000000000000000";
    input_dim2x_x1_at_entry_1992 <= "0000000000000000";
    ptr_deref_2100_word_offset_0 <= "00000000000000";
    ptr_deref_2125_word_offset_0 <= "00000000000000";
    type_cast_1903_wire_constant <= "00000000000000000000000000010000";
    type_cast_1931_wire_constant <= "0000000000000010";
    type_cast_1937_wire_constant <= "1111111111111111";
    type_cast_1948_wire_constant <= "1111111111111111";
    type_cast_1967_wire_constant <= "1111111111111100";
    type_cast_1982_wire_constant <= "00000000000000000000000000000001";
    type_cast_2105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2111_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2145_wire_constant <= "0000000000000100";
    type_cast_2155_wire_constant <= "0000000000000000";
    type_cast_2165_wire_constant <= "0000000000000001";
    type_cast_2196_wire_constant <= "0000000000000000";
    type_cast_2212_wire_constant <= "00000000000000000000000000000001";
    type_cast_2229_wire_constant <= "0000000000000001";
    phi_stmt_2002: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2005_wire;
      req(0) <= phi_stmt_2002_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2002",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2002_ack_0,
          idata => idata,
          odata => input_dim0x_x1_at_entry_2002,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2002
    phi_stmt_2009: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2012_wire & indvar_at_entry_1987;
      req <= phi_stmt_2009_req_0 & phi_stmt_2009_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2009",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2009_ack_0,
          idata => idata,
          odata => indvar_2009,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2009
    phi_stmt_2014: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim2x_x1_at_entry_1992 & type_cast_2018_wire;
      req <= phi_stmt_2014_req_0 & phi_stmt_2014_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2014",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2014_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2014,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2014
    phi_stmt_2019: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim1x_x1_at_entry_1997 & type_cast_2023_wire;
      req <= phi_stmt_2019_req_0 & phi_stmt_2019_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2019",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2019_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2019,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2019
    phi_stmt_2024: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2027_wire & input_dim0x_x1_at_entry_2002_2028_buffered;
      req <= phi_stmt_2024_req_0 & phi_stmt_2024_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2024",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2024_ack_0,
          idata => idata,
          odata => input_dim0x_x1_2024,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2024
    -- flow-through select operator MUX_2156_inst
    input_dim2x_x0_2157 <= add101_2129_delayed_1_0_2150 when (cmp_2141(0) /=  '0') else type_cast_2155_wire_constant;
    -- flow-through select operator MUX_2198_inst
    input_dim1x_x2_2199 <= type_cast_2196_wire_constant when (cmp109_2180(0) /=  '0') else input_dim1x_x0_2175;
    W_add101_2129_delayed_1_0_2148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add101_2129_delayed_1_0_2148_inst_req_0;
      W_add101_2129_delayed_1_0_2148_inst_ack_0<= wack(0);
      rreq(0) <= W_add101_2129_delayed_1_0_2148_inst_req_1;
      W_add101_2129_delayed_1_0_2148_inst_ack_1<= rack(0);
      W_add101_2129_delayed_1_0_2148_inst : InterlockBuffer generic map ( -- 
        name => "W_add101_2129_delayed_1_0_2148_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add101_2147,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add101_2129_delayed_1_0_2150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx86_2106_delayed_6_0_2121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx86_2106_delayed_6_0_2121_inst_req_0;
      W_arrayidx86_2106_delayed_6_0_2121_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx86_2106_delayed_6_0_2121_inst_req_1;
      W_arrayidx86_2106_delayed_6_0_2121_inst_ack_1<= rack(0);
      W_arrayidx86_2106_delayed_6_0_2121_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx86_2106_delayed_6_0_2121_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx86_2120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_2106_delayed_6_0_2123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim0x_x1_2160_delayed_3_0_2185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim0x_x1_2160_delayed_3_0_2185_inst_req_0;
      W_input_dim0x_x1_2160_delayed_3_0_2185_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim0x_x1_2160_delayed_3_0_2185_inst_req_1;
      W_input_dim0x_x1_2160_delayed_3_0_2185_inst_ack_1<= rack(0);
      W_input_dim0x_x1_2160_delayed_3_0_2185_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim0x_x1_2160_delayed_3_0_2185_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_2024,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_2160_delayed_3_0_2187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim1x_x1_2146_delayed_2_0_2168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim1x_x1_2146_delayed_2_0_2168_inst_req_0;
      W_input_dim1x_x1_2146_delayed_2_0_2168_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim1x_x1_2146_delayed_2_0_2168_inst_req_1;
      W_input_dim1x_x1_2146_delayed_2_0_2168_inst_ack_1<= rack(0);
      W_input_dim1x_x1_2146_delayed_2_0_2168_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim1x_x1_2146_delayed_2_0_2168_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2019,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim1x_x1_2146_delayed_2_0_2170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_2215_inst
    process(cmp121_2208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp121_2208(0 downto 0);
      whilex_xbody_whilex_xend_taken_2217 <= tmp_var; -- 
    end process;
    addr_of_2096_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2096_final_reg_req_0;
      addr_of_2096_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2096_final_reg_req_1;
      addr_of_2096_final_reg_ack_1<= rack(0);
      addr_of_2096_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2096_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2095_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx81_2097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2119_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2119_final_reg_req_0;
      addr_of_2119_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2119_final_reg_req_1;
      addr_of_2119_final_reg_ack_1<= rack(0);
      addr_of_2119_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2119_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2118_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_2120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    input_dim0x_x1_at_entry_2002_2028_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= input_dim0x_x1_at_entry_2002_2028_buf_req_0;
      input_dim0x_x1_at_entry_2002_2028_buf_ack_0<= wack(0);
      rreq(0) <= input_dim0x_x1_at_entry_2002_2028_buf_req_1;
      input_dim0x_x1_at_entry_2002_2028_buf_ack_1<= rack(0);
      input_dim0x_x1_at_entry_2002_2028_buf : InterlockBuffer generic map ( -- 
        name => "input_dim0x_x1_at_entry_2002_2028_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_at_entry_2002,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_at_entry_2002_2028_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1898_inst_req_0;
      type_cast_1898_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1898_inst_req_1;
      type_cast_1898_inst_ack_1<= rack(0);
      type_cast_1898_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1898_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1911_inst_req_0;
      type_cast_1911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1911_inst_req_1;
      type_cast_1911_inst_ack_1<= rack(0);
      type_cast_1911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1912,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1958_inst_req_0;
      type_cast_1958_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1958_inst_req_1;
      type_cast_1958_inst_ack_1<= rack(0);
      type_cast_1958_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1959,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1962_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1962_inst_req_0;
      type_cast_1962_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1962_inst_req_1;
      type_cast_1962_inst_ack_1<= rack(0);
      type_cast_1962_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1962_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1923,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1973_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1973_inst_req_0;
      type_cast_1973_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1973_inst_req_1;
      type_cast_1973_inst_ack_1<= rack(0);
      type_cast_1973_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1973_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1972_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_1974,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1977_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1977_inst_req_0;
      type_cast_1977_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1977_inst_req_1;
      type_cast_1977_inst_ack_1<= rack(0);
      type_cast_1977_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1977_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_1978,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2005_inst_req_0;
      type_cast_2005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2005_inst_req_1;
      type_cast_2005_inst_ack_1<= rack(0);
      type_cast_2005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr134_1933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2005_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2012_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2012_inst_req_0;
      type_cast_2012_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2012_inst_req_1;
      type_cast_2012_inst_ack_1<= rack(0);
      type_cast_2012_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2012_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2012_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2018_inst_req_0;
      type_cast_2018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2018_inst_req_1;
      type_cast_2018_inst_ack_1<= rack(0);
      type_cast_2018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2018_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0_2157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2018_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2023_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2023_inst_req_0;
      type_cast_2023_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2023_inst_req_1;
      type_cast_2023_inst_ack_1<= rack(0);
      type_cast_2023_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2023_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2023_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2027_inst_req_0;
      type_cast_2027_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2027_inst_req_1;
      type_cast_2027_inst_ack_1<= rack(0);
      type_cast_2027_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2027_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc113x_xinput_dim0x_x1_2192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2027_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2057_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2057_inst_req_0;
      type_cast_2057_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2057_inst_req_1;
      type_cast_2057_inst_ack_1<= rack(0);
      type_cast_2057_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2057_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2014,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2058,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2061_inst_req_0;
      type_cast_2061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2061_inst_req_1;
      type_cast_2061_inst_ack_1<= rack(0);
      type_cast_2061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2054,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2065_inst_req_0;
      type_cast_2065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2065_inst_req_1;
      type_cast_2065_inst_ack_1<= rack(0);
      type_cast_2065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2044,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2066,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2089_inst_req_0;
      type_cast_2089_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2089_inst_req_1;
      type_cast_2089_inst_ack_1<= rack(0);
      type_cast_2089_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_src_0x_x0_2034,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2090,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2130_inst_req_0;
      type_cast_2130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2130_inst_req_1;
      type_cast_2130_inst_ack_1<= rack(0);
      type_cast_2130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2130_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2014,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2134_inst_req_0;
      type_cast_2134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2134_inst_req_1;
      type_cast_2134_inst_ack_1<= rack(0);
      type_cast_2134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2134_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv97_1974,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2118_2118_delayed_2_0_2135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2138_inst
    process(conv95_2131) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv95_2131(31 downto 0);
      type_cast_2138_wire <= tmp_var; -- 
    end process;
    type_cast_2160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2160_inst_req_0;
      type_cast_2160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2160_inst_req_1;
      type_cast_2160_inst_ack_1<= rack(0);
      type_cast_2160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2160_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_2141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_18_2161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2183_inst_req_0;
      type_cast_2183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2183_inst_req_1;
      type_cast_2183_inst_ack_1<= rack(0);
      type_cast_2183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2183_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp109_2180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc113_2184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2202_inst_req_0;
      type_cast_2202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2202_inst_req_1;
      type_cast_2202_inst_ack_1<= rack(0);
      type_cast_2202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc113x_xinput_dim0x_x1_2192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_2203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2095_index_1_rename
    process(R_idxprom_2094_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2094_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2094_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2095_index_1_resize
    process(idxprom_2090) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2090;
      ov := iv(13 downto 0);
      R_idxprom_2094_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2095_root_address_inst
    process(array_obj_ref_2095_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2095_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2095_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2118_index_1_rename
    process(R_idxprom85_2117_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom85_2117_resized;
      ov(13 downto 0) := iv;
      R_idxprom85_2117_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2118_index_1_resize
    process(idxprom85_2113) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom85_2113;
      ov := iv(13 downto 0);
      R_idxprom85_2117_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2118_root_address_inst
    process(array_obj_ref_2118_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2118_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2118_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_addr_0
    process(ptr_deref_2100_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2100_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_base_resize
    process(arrayidx81_2097) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx81_2097;
      ov := iv(13 downto 0);
      ptr_deref_2100_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_gather_scatter
    process(ptr_deref_2100_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_data_0;
      ov(63 downto 0) := iv;
      tmp82_2101 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_root_address_inst
    process(ptr_deref_2100_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2100_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2125_addr_0
    process(ptr_deref_2125_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2125_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2125_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2125_base_resize
    process(arrayidx86_2106_delayed_6_0_2123) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx86_2106_delayed_6_0_2123;
      ov := iv(13 downto 0);
      ptr_deref_2125_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2125_gather_scatter
    process(tmp82_2101) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp82_2101;
      ov(63 downto 0) := iv;
      ptr_deref_2125_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2125_root_address_inst
    process(ptr_deref_2125_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2125_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2125_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_2007_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2220_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2007_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2007_branch_req_0,
          ack0 => do_while_stmt_2007_branch_ack_0,
          ack1 => do_while_stmt_2007_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2221_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_2217;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2221_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2221_branch_req_0,
          ack0 => if_stmt_2221_branch_ack_0,
          ack1 => if_stmt_2221_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1938_inst
    process(call7_1880) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1880, type_cast_1937_wire_constant, tmp_var);
      add45_1939 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1949_inst
    process(call9_1883) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1883, type_cast_1948_wire_constant, tmp_var);
      add58_1950 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1968_inst
    process(call3_1874) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call3_1874, type_cast_1967_wire_constant, tmp_var);
      sub91_1969 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2043_inst
    process(sub_1944, mul_2039) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1944, mul_2039, tmp_var);
      sub48_2044 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2053_inst
    process(sub61_1955, mul54_2049) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1955, mul54_2049, tmp_var);
      sub62_2054 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2146_inst
    process(input_dim2x_x1_2014) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2014, type_cast_2145_wire_constant, tmp_var);
      add101_2147 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2174_inst
    process(inc_2167, input_dim1x_x1_2146_delayed_2_0_2170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc_2167, input_dim1x_x1_2146_delayed_2_0_2170, tmp_var);
      input_dim1x_x0_2175 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2191_inst
    process(inc113_2184, input_dim0x_x1_2160_delayed_3_0_2187) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc113_2184, input_dim0x_x1_2160_delayed_3_0_2187, tmp_var);
      inc113x_xinput_dim0x_x1_2192 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2033_inst
    process(add_1917, indvar_2009) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1917, indvar_2009, tmp_var);
      add_src_0x_x0_2034 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2213_inst
    process(indvar_2009) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2009, type_cast_2212_wire_constant, tmp_var);
      indvarx_xnext_2214 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2075_inst
    process(mul76_2071, conv70_2062) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2071, conv70_2062, tmp_var);
      add77_2076 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2085_inst
    process(mul78_2081, conv65_2058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2081, conv65_2058, tmp_var);
      add79_2086 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2112_inst
    process(shr84_2107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr84_2107, type_cast_2111_wire_constant, tmp_var);
      idxprom85_2113 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2179_inst
    process(input_dim1x_x0_2175, call1_1871) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1x_x0_2175, call1_1871, tmp_var);
      cmp109_2180 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2207_inst
    process(conv116_2203, shr120135_1984) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv116_2203, shr120135_1984, tmp_var);
      cmp121_2208 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1932_inst
    process(call_1868) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1868, type_cast_1931_wire_constant, tmp_var);
      shr134_1933 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1983_inst
    process(conv119_1978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv119_1978, type_cast_1982_wire_constant, tmp_var);
      shr120135_1984 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2106_inst
    process(add79_2086) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2086, type_cast_2105_wire_constant, tmp_var);
      shr84_2107 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2038_inst
    process(input_dim0x_x1_2024, call13_1889) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x1_2024, call13_1889, tmp_var);
      mul_2039 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2048_inst
    process(input_dim1x_x1_2019, call13_1889) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2019, call13_1889, tmp_var);
      mul54_2049 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2070_inst
    process(conv75_2066, conv73_1963) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2066, conv73_1963, tmp_var);
      mul76_2071 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2080_inst
    process(add77_2076, conv68_1959) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2076, conv68_1959, tmp_var);
      mul78_2081 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2220_inst
    process(cmp121_2208) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp121_2208, tmp_var);
      NOT_u1_u1_2220_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u32_u32_1916_inst
    process(shl_1905, conv17_1912) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1905, conv17_1912, tmp_var);
      add_1917 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1904_inst
    process(conv_1899) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1899, type_cast_1903_wire_constant, tmp_var);
      shl_1905 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2140_inst
    process(type_cast_2138_wire, type_cast_2118_2118_delayed_2_0_2135) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2138_wire, type_cast_2118_2118_delayed_2_0_2135, tmp_var);
      cmp_2141 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1943_inst
    process(add45_1939, call14_1892) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1939, call14_1892, tmp_var);
      sub_1944 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1954_inst
    process(add58_1950, call14_1892) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1950, call14_1892, tmp_var);
      sub61_1955 <= tmp_var; --
    end process;
    -- binary operator XOR_u16_u16_2166_inst
    process(iNsTr_18_2161) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntXor_proc(iNsTr_18_2161, type_cast_2165_wire_constant, tmp_var);
      inc_2167 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2095_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2094_scaled;
      array_obj_ref_2095_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2095_index_offset_req_0;
      array_obj_ref_2095_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2095_index_offset_req_1;
      array_obj_ref_2095_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2118_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom85_2117_scaled;
      array_obj_ref_2118_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2118_index_offset_req_0;
      array_obj_ref_2118_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2118_index_offset_req_1;
      array_obj_ref_2118_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- unary operator type_cast_1972_inst
    process(sub91_1969) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", sub91_1969, tmp_var);
      type_cast_1972_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2100_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2100_load_0_req_0;
      ptr_deref_2100_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2100_load_0_req_1;
      ptr_deref_2100_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2100_word_address_0;
      ptr_deref_2100_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2125_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2125_store_0_req_0;
      ptr_deref_2125_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2125_store_0_req_1;
      ptr_deref_2125_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2125_word_address_0;
      data_in <= ptr_deref_2125_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1907_inst RPIPE_Block1_start_1925_inst RPIPE_Block1_start_1922_inst RPIPE_Block1_start_1894_inst RPIPE_Block1_start_1876_inst RPIPE_Block1_start_1891_inst RPIPE_Block1_start_1888_inst RPIPE_Block1_start_1919_inst RPIPE_Block1_start_1885_inst RPIPE_Block1_start_1873_inst RPIPE_Block1_start_1882_inst RPIPE_Block1_start_1870_inst RPIPE_Block1_start_1867_inst RPIPE_Block1_start_1879_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1907_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1925_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1922_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1894_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1876_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1891_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1888_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1919_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1885_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1873_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1882_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1870_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1867_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1879_inst_req_0;
      RPIPE_Block1_start_1907_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1925_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1922_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1894_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1876_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1891_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1888_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1919_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1885_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1873_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1882_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1870_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1867_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1879_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1907_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1925_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1922_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1894_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1876_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1891_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1888_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1919_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1885_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1873_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1882_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1870_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1867_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1879_inst_req_1;
      RPIPE_Block1_start_1907_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1925_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1922_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1894_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1876_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1891_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1888_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1919_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1885_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1873_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1882_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1870_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1867_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1879_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call16_1908 <= data_out(223 downto 208);
      call22_1926 <= data_out(207 downto 192);
      call20_1923 <= data_out(191 downto 176);
      call15_1895 <= data_out(175 downto 160);
      call5_1877 <= data_out(159 downto 144);
      call14_1892 <= data_out(143 downto 128);
      call13_1889 <= data_out(127 downto 112);
      call18_1920 <= data_out(111 downto 96);
      call11_1886 <= data_out(95 downto 80);
      call3_1874 <= data_out(79 downto 64);
      call9_1883 <= data_out(63 downto 48);
      call1_1871 <= data_out(47 downto 32);
      call_1868 <= data_out(31 downto 16);
      call7_1880 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2227_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2227_inst_req_0;
      WPIPE_Block1_done_2227_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2227_inst_req_1;
      WPIPE_Block1_done_2227_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2229_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5701_start: Boolean;
  signal convTransposeC_CP_5701_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2394_inst_ack_1 : boolean;
  signal type_cast_2439_inst_ack_0 : boolean;
  signal do_while_stmt_2389_branch_req_0 : boolean;
  signal phi_stmt_2396_req_0 : boolean;
  signal type_cast_2333_inst_req_1 : boolean;
  signal phi_stmt_2396_ack_0 : boolean;
  signal type_cast_2439_inst_req_0 : boolean;
  signal type_cast_2344_inst_req_1 : boolean;
  signal phi_stmt_2401_ack_0 : boolean;
  signal RPIPE_Block2_start_2296_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2293_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2290_inst_ack_1 : boolean;
  signal type_cast_2404_inst_ack_1 : boolean;
  signal type_cast_2282_inst_req_1 : boolean;
  signal type_cast_2344_inst_ack_1 : boolean;
  signal type_cast_2394_inst_req_1 : boolean;
  signal type_cast_2348_inst_req_1 : boolean;
  signal type_cast_2394_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2293_inst_ack_0 : boolean;
  signal type_cast_2269_inst_ack_1 : boolean;
  signal type_cast_2443_inst_ack_1 : boolean;
  signal type_cast_2439_inst_ack_1 : boolean;
  signal input_dim0x_x1_at_entry_2384_2410_buf_req_0 : boolean;
  signal type_cast_2439_inst_req_1 : boolean;
  signal type_cast_2282_inst_req_0 : boolean;
  signal type_cast_2443_inst_req_0 : boolean;
  signal type_cast_2443_inst_ack_0 : boolean;
  signal type_cast_2443_inst_req_1 : boolean;
  signal type_cast_2409_inst_req_0 : boolean;
  signal type_cast_2333_inst_ack_1 : boolean;
  signal phi_stmt_2401_req_0 : boolean;
  signal phi_stmt_2406_ack_0 : boolean;
  signal phi_stmt_2406_req_0 : boolean;
  signal type_cast_2394_inst_ack_0 : boolean;
  signal phi_stmt_2406_req_1 : boolean;
  signal type_cast_2282_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2278_inst_req_0 : boolean;
  signal type_cast_2404_inst_req_1 : boolean;
  signal type_cast_2344_inst_ack_0 : boolean;
  signal type_cast_2269_inst_req_1 : boolean;
  signal type_cast_2409_inst_ack_0 : boolean;
  signal type_cast_2348_inst_ack_0 : boolean;
  signal phi_stmt_2396_req_1 : boolean;
  signal input_dim0x_x1_at_entry_2384_2410_buf_ack_1 : boolean;
  signal type_cast_2348_inst_req_0 : boolean;
  signal type_cast_2409_inst_req_1 : boolean;
  signal type_cast_2404_inst_ack_0 : boolean;
  signal type_cast_2447_inst_req_0 : boolean;
  signal type_cast_2447_inst_ack_0 : boolean;
  signal type_cast_2404_inst_req_0 : boolean;
  signal type_cast_2409_inst_ack_1 : boolean;
  signal input_dim0x_x1_at_entry_2384_2410_buf_ack_0 : boolean;
  signal type_cast_2447_inst_req_1 : boolean;
  signal type_cast_2447_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2278_inst_ack_1 : boolean;
  signal input_dim0x_x1_at_entry_2384_2410_buf_req_1 : boolean;
  signal RPIPE_Block2_start_2278_inst_req_1 : boolean;
  signal type_cast_2344_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2296_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2290_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2238_inst_req_0 : boolean;
  signal type_cast_2333_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_req_1 : boolean;
  signal type_cast_2333_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2238_inst_ack_1 : boolean;
  signal phi_stmt_2401_req_1 : boolean;
  signal RPIPE_Block2_start_2241_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2241_inst_ack_0 : boolean;
  signal type_cast_2399_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2241_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2241_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2296_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2296_inst_req_0 : boolean;
  signal type_cast_2399_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2244_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2244_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2244_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2244_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2290_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2278_inst_ack_0 : boolean;
  signal type_cast_2348_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2247_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2247_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2290_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2247_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2247_inst_ack_1 : boolean;
  signal phi_stmt_2391_ack_0 : boolean;
  signal type_cast_2399_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2250_inst_req_0 : boolean;
  signal type_cast_2329_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2250_inst_ack_0 : boolean;
  signal type_cast_2399_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2250_inst_req_1 : boolean;
  signal type_cast_2329_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2250_inst_ack_1 : boolean;
  signal phi_stmt_2391_req_1 : boolean;
  signal RPIPE_Block2_start_2293_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2253_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2253_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2253_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2253_inst_ack_1 : boolean;
  signal phi_stmt_2391_req_0 : boolean;
  signal RPIPE_Block2_start_2293_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2256_inst_req_0 : boolean;
  signal type_cast_2329_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2256_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2256_inst_req_1 : boolean;
  signal type_cast_2329_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2256_inst_ack_1 : boolean;
  signal type_cast_2282_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2259_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2259_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2259_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2259_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2262_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2262_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2262_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2262_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2265_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2265_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2265_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2265_inst_ack_1 : boolean;
  signal type_cast_2269_inst_req_0 : boolean;
  signal type_cast_2269_inst_ack_0 : boolean;
  signal type_cast_2471_inst_req_0 : boolean;
  signal type_cast_2471_inst_ack_0 : boolean;
  signal type_cast_2471_inst_req_1 : boolean;
  signal type_cast_2471_inst_ack_1 : boolean;
  signal array_obj_ref_2477_index_offset_req_0 : boolean;
  signal array_obj_ref_2477_index_offset_ack_0 : boolean;
  signal array_obj_ref_2477_index_offset_req_1 : boolean;
  signal array_obj_ref_2477_index_offset_ack_1 : boolean;
  signal addr_of_2478_final_reg_req_0 : boolean;
  signal addr_of_2478_final_reg_ack_0 : boolean;
  signal addr_of_2478_final_reg_req_1 : boolean;
  signal addr_of_2478_final_reg_ack_1 : boolean;
  signal ptr_deref_2482_load_0_req_0 : boolean;
  signal ptr_deref_2482_load_0_ack_0 : boolean;
  signal ptr_deref_2482_load_0_req_1 : boolean;
  signal ptr_deref_2482_load_0_ack_1 : boolean;
  signal array_obj_ref_2500_index_offset_req_0 : boolean;
  signal array_obj_ref_2500_index_offset_ack_0 : boolean;
  signal array_obj_ref_2500_index_offset_req_1 : boolean;
  signal array_obj_ref_2500_index_offset_ack_1 : boolean;
  signal addr_of_2501_final_reg_req_0 : boolean;
  signal addr_of_2501_final_reg_ack_0 : boolean;
  signal addr_of_2501_final_reg_req_1 : boolean;
  signal addr_of_2501_final_reg_ack_1 : boolean;
  signal W_arrayidx86_2473_delayed_6_0_2503_inst_req_0 : boolean;
  signal W_arrayidx86_2473_delayed_6_0_2503_inst_ack_0 : boolean;
  signal W_arrayidx86_2473_delayed_6_0_2503_inst_req_1 : boolean;
  signal W_arrayidx86_2473_delayed_6_0_2503_inst_ack_1 : boolean;
  signal ptr_deref_2507_store_0_req_0 : boolean;
  signal ptr_deref_2507_store_0_ack_0 : boolean;
  signal ptr_deref_2507_store_0_req_1 : boolean;
  signal ptr_deref_2507_store_0_ack_1 : boolean;
  signal type_cast_2512_inst_req_0 : boolean;
  signal type_cast_2512_inst_ack_0 : boolean;
  signal type_cast_2512_inst_req_1 : boolean;
  signal type_cast_2512_inst_ack_1 : boolean;
  signal type_cast_2516_inst_req_0 : boolean;
  signal type_cast_2516_inst_ack_0 : boolean;
  signal type_cast_2516_inst_req_1 : boolean;
  signal type_cast_2516_inst_ack_1 : boolean;
  signal W_add101_2496_delayed_1_0_2530_inst_req_0 : boolean;
  signal W_add101_2496_delayed_1_0_2530_inst_ack_0 : boolean;
  signal W_add101_2496_delayed_1_0_2530_inst_req_1 : boolean;
  signal W_add101_2496_delayed_1_0_2530_inst_ack_1 : boolean;
  signal type_cast_2542_inst_req_0 : boolean;
  signal type_cast_2542_inst_ack_0 : boolean;
  signal type_cast_2542_inst_req_1 : boolean;
  signal type_cast_2542_inst_ack_1 : boolean;
  signal W_input_dim1x_x1_2513_delayed_2_0_2550_inst_req_0 : boolean;
  signal W_input_dim1x_x1_2513_delayed_2_0_2550_inst_ack_0 : boolean;
  signal W_input_dim1x_x1_2513_delayed_2_0_2550_inst_req_1 : boolean;
  signal W_input_dim1x_x1_2513_delayed_2_0_2550_inst_ack_1 : boolean;
  signal type_cast_2565_inst_req_0 : boolean;
  signal type_cast_2565_inst_ack_0 : boolean;
  signal type_cast_2565_inst_req_1 : boolean;
  signal type_cast_2565_inst_ack_1 : boolean;
  signal W_input_dim0x_x1_2527_delayed_3_0_2567_inst_req_0 : boolean;
  signal W_input_dim0x_x1_2527_delayed_3_0_2567_inst_ack_0 : boolean;
  signal W_input_dim0x_x1_2527_delayed_3_0_2567_inst_req_1 : boolean;
  signal W_input_dim0x_x1_2527_delayed_3_0_2567_inst_ack_1 : boolean;
  signal type_cast_2584_inst_req_0 : boolean;
  signal type_cast_2584_inst_ack_0 : boolean;
  signal type_cast_2584_inst_req_1 : boolean;
  signal type_cast_2584_inst_ack_1 : boolean;
  signal do_while_stmt_2389_branch_ack_0 : boolean;
  signal do_while_stmt_2389_branch_ack_1 : boolean;
  signal if_stmt_2603_branch_req_0 : boolean;
  signal if_stmt_2603_branch_ack_1 : boolean;
  signal if_stmt_2603_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2609_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2609_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2609_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2609_inst_ack_1 : boolean;
  signal type_cast_2387_inst_req_0 : boolean;
  signal type_cast_2387_inst_ack_0 : boolean;
  signal type_cast_2387_inst_req_1 : boolean;
  signal type_cast_2387_inst_ack_1 : boolean;
  signal phi_stmt_2384_req_0 : boolean;
  signal phi_stmt_2384_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5701_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5701_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5701_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5701_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5701: Block -- control-path 
    signal convTransposeC_CP_5701_elements: BooleanArray(226 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5701_elements(0) <= convTransposeC_CP_5701_start;
    convTransposeC_CP_5701_symbol <= convTransposeC_CP_5701_elements(222);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2236/$entry
      -- CP-element group 0: 	 branch_block_stmt_2236/branch_block_stmt_2236__entry__
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297__entry__
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/$entry
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_update_start_
      -- 
    cr_5908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(0), ack => type_cast_2282_inst_req_1); -- 
    cr_5880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(0), ack => type_cast_2269_inst_req_1); -- 
    rr_5735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(0), ack => RPIPE_Block2_start_2238_inst_req_0); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	218 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	219 
    -- CP-element group 1: 	220 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_2236/do_while_stmt_2389__exit__
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603__entry__
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_2236/R_whilex_xbody_whilex_xend_taken_2604_place
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_2236/if_stmt_2603_else_link/$entry
      -- 
    branch_req_6608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(1), ack => if_stmt_2603_branch_req_0); -- 
    convTransposeC_CP_5701_elements(1) <= convTransposeC_CP_5701_elements(218);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Update/cr
      -- 
    ra_5736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2238_inst_ack_0, ack => convTransposeC_CP_5701_elements(2)); -- 
    cr_5740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(2), ack => RPIPE_Block2_start_2238_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2238_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Sample/rr
      -- 
    ca_5741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2238_inst_ack_1, ack => convTransposeC_CP_5701_elements(3)); -- 
    rr_5749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(3), ack => RPIPE_Block2_start_2241_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Update/cr
      -- 
    ra_5750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2241_inst_ack_0, ack => convTransposeC_CP_5701_elements(4)); -- 
    cr_5754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(4), ack => RPIPE_Block2_start_2241_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2241_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Sample/rr
      -- 
    ca_5755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2241_inst_ack_1, ack => convTransposeC_CP_5701_elements(5)); -- 
    rr_5763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(5), ack => RPIPE_Block2_start_2244_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Update/cr
      -- 
    ra_5764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2244_inst_ack_0, ack => convTransposeC_CP_5701_elements(6)); -- 
    cr_5768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(6), ack => RPIPE_Block2_start_2244_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2244_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Sample/rr
      -- 
    ca_5769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2244_inst_ack_1, ack => convTransposeC_CP_5701_elements(7)); -- 
    rr_5777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(7), ack => RPIPE_Block2_start_2247_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Update/cr
      -- 
    ra_5778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2247_inst_ack_0, ack => convTransposeC_CP_5701_elements(8)); -- 
    cr_5782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(8), ack => RPIPE_Block2_start_2247_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2247_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Sample/rr
      -- 
    ca_5783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2247_inst_ack_1, ack => convTransposeC_CP_5701_elements(9)); -- 
    rr_5791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(9), ack => RPIPE_Block2_start_2250_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Update/cr
      -- 
    ra_5792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2250_inst_ack_0, ack => convTransposeC_CP_5701_elements(10)); -- 
    cr_5796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(10), ack => RPIPE_Block2_start_2250_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2250_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Sample/rr
      -- 
    ca_5797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2250_inst_ack_1, ack => convTransposeC_CP_5701_elements(11)); -- 
    rr_5805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(11), ack => RPIPE_Block2_start_2253_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Update/cr
      -- 
    ra_5806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2253_inst_ack_0, ack => convTransposeC_CP_5701_elements(12)); -- 
    cr_5810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(12), ack => RPIPE_Block2_start_2253_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2253_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Sample/rr
      -- 
    ca_5811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2253_inst_ack_1, ack => convTransposeC_CP_5701_elements(13)); -- 
    rr_5819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(13), ack => RPIPE_Block2_start_2256_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Update/cr
      -- 
    ra_5820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2256_inst_ack_0, ack => convTransposeC_CP_5701_elements(14)); -- 
    cr_5824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(14), ack => RPIPE_Block2_start_2256_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2256_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Sample/rr
      -- 
    ca_5825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2256_inst_ack_1, ack => convTransposeC_CP_5701_elements(15)); -- 
    rr_5833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(15), ack => RPIPE_Block2_start_2259_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Update/cr
      -- 
    ra_5834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2259_inst_ack_0, ack => convTransposeC_CP_5701_elements(16)); -- 
    cr_5838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(16), ack => RPIPE_Block2_start_2259_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2259_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Sample/rr
      -- 
    ca_5839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2259_inst_ack_1, ack => convTransposeC_CP_5701_elements(17)); -- 
    rr_5847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(17), ack => RPIPE_Block2_start_2262_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Update/cr
      -- 
    ra_5848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2262_inst_ack_0, ack => convTransposeC_CP_5701_elements(18)); -- 
    cr_5852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(18), ack => RPIPE_Block2_start_2262_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2262_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Sample/rr
      -- 
    ca_5853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2262_inst_ack_1, ack => convTransposeC_CP_5701_elements(19)); -- 
    rr_5861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(19), ack => RPIPE_Block2_start_2265_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Update/cr
      -- 
    ra_5862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2265_inst_ack_0, ack => convTransposeC_CP_5701_elements(20)); -- 
    cr_5866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(20), ack => RPIPE_Block2_start_2265_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2265_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Sample/rr
      -- 
    ca_5867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2265_inst_ack_1, ack => convTransposeC_CP_5701_elements(21)); -- 
    rr_5875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(21), ack => type_cast_2269_inst_req_0); -- 
    rr_5889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(21), ack => RPIPE_Block2_start_2278_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Sample/ra
      -- 
    ra_5876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_0, ack => convTransposeC_CP_5701_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2269_update_completed_
      -- 
    ca_5881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2269_inst_ack_1, ack => convTransposeC_CP_5701_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Sample/ra
      -- 
    ra_5890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2278_inst_ack_0, ack => convTransposeC_CP_5701_elements(24)); -- 
    cr_5894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(24), ack => RPIPE_Block2_start_2278_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2278_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_sample_start_
      -- 
    ca_5895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2278_inst_ack_1, ack => convTransposeC_CP_5701_elements(25)); -- 
    rr_5903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(25), ack => type_cast_2282_inst_req_0); -- 
    rr_5917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(25), ack => RPIPE_Block2_start_2290_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_sample_completed_
      -- 
    ra_5904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_0, ack => convTransposeC_CP_5701_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/type_cast_2282_Update/ca
      -- 
    ca_5909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_1, ack => convTransposeC_CP_5701_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_sample_completed_
      -- 
    ra_5918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2290_inst_ack_0, ack => convTransposeC_CP_5701_elements(28)); -- 
    cr_5922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(28), ack => RPIPE_Block2_start_2290_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2290_update_completed_
      -- 
    ca_5923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2290_inst_ack_1, ack => convTransposeC_CP_5701_elements(29)); -- 
    rr_5931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(29), ack => RPIPE_Block2_start_2293_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Update/$entry
      -- 
    ra_5932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2293_inst_ack_0, ack => convTransposeC_CP_5701_elements(30)); -- 
    cr_5936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(30), ack => RPIPE_Block2_start_2293_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2293_Update/$exit
      -- 
    ca_5937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2293_inst_ack_1, ack => convTransposeC_CP_5701_elements(31)); -- 
    rr_5945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(31), ack => RPIPE_Block2_start_2296_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_sample_completed_
      -- 
    ra_5946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2296_inst_ack_0, ack => convTransposeC_CP_5701_elements(32)); -- 
    cr_5950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(32), ack => RPIPE_Block2_start_2296_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/RPIPE_Block2_start_2296_update_completed_
      -- 
    ca_5951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2296_inst_ack_1, ack => convTransposeC_CP_5701_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297__exit__
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366__entry__
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2239_to_assign_stmt_2297/$exit
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Sample/rr
      -- 
    cr_5981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2333_inst_req_1); -- 
    cr_5995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2344_inst_req_1); -- 
    cr_6009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2348_inst_req_1); -- 
    rr_6004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2348_inst_req_0); -- 
    rr_5990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2344_inst_req_0); -- 
    rr_5976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2333_inst_req_0); -- 
    cr_5967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2329_inst_req_1); -- 
    rr_5962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(34), ack => type_cast_2329_inst_req_0); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(23) & convTransposeC_CP_5701_elements(27) & convTransposeC_CP_5701_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Sample/ra
      -- 
    ra_5963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2329_inst_ack_0, ack => convTransposeC_CP_5701_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2329_Update/$exit
      -- 
    ca_5968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2329_inst_ack_1, ack => convTransposeC_CP_5701_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_sample_completed_
      -- 
    ra_5977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2333_inst_ack_0, ack => convTransposeC_CP_5701_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2333_update_completed_
      -- 
    ca_5982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2333_inst_ack_1, ack => convTransposeC_CP_5701_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Sample/$exit
      -- 
    ra_5991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2344_inst_ack_0, ack => convTransposeC_CP_5701_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2344_update_completed_
      -- 
    ca_5996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2344_inst_ack_1, ack => convTransposeC_CP_5701_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_sample_completed_
      -- 
    ra_6005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2348_inst_ack_0, ack => convTransposeC_CP_5701_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/type_cast_2348_Update/ca
      -- 
    ca_6010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2348_inst_ack_1, ack => convTransposeC_CP_5701_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	223 
    -- CP-element group 43: 	224 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366/$exit
      -- CP-element group 43: 	 branch_block_stmt_2236/assign_stmt_2304_to_assign_stmt_2366__exit__
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Update/cr
      -- 
    rr_6654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(43), ack => type_cast_2387_inst_req_0); -- 
    cr_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(43), ack => type_cast_2387_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(36) & convTransposeC_CP_5701_elements(38) & convTransposeC_CP_5701_elements(40) & convTransposeC_CP_5701_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	226 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	50 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_2236/do_while_stmt_2389/$entry
      -- CP-element group 44: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389__entry__
      -- 
    convTransposeC_CP_5701_elements(44) <= convTransposeC_CP_5701_elements(226);
    -- CP-element group 45:  merge  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	218 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389__exit__
      -- 
    -- Element group convTransposeC_CP_5701_elements(45) is bound as output of CP function.
    -- CP-element group 46:  merge  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_back
      -- 
    -- Element group convTransposeC_CP_5701_elements(46) is bound as output of CP function.
    -- CP-element group 47:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	52 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	217 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2236/do_while_stmt_2389/condition_done
      -- CP-element group 47: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_exit/$entry
      -- CP-element group 47: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_taken/$entry
      -- 
    convTransposeC_CP_5701_elements(47) <= convTransposeC_CP_5701_elements(52);
    -- CP-element group 48:  branch  place  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	215 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_body_done
      -- 
    convTransposeC_CP_5701_elements(48) <= convTransposeC_CP_5701_elements(215);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	61 
    -- CP-element group 49: 	82 
    -- CP-element group 49: 	103 
    -- CP-element group 49: 	124 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/back_edge_to_loop_body
      -- 
    convTransposeC_CP_5701_elements(49) <= convTransposeC_CP_5701_elements(46);
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	44 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	63 
    -- CP-element group 50: 	84 
    -- CP-element group 50: 	105 
    -- CP-element group 50: 	126 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/first_time_through_loop_body
      -- 
    convTransposeC_CP_5701_elements(50) <= convTransposeC_CP_5701_elements(44);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	57 
    -- CP-element group 51: 	58 
    -- CP-element group 51: 	76 
    -- CP-element group 51: 	77 
    -- CP-element group 51: 	97 
    -- CP-element group 51: 	98 
    -- CP-element group 51: 	118 
    -- CP-element group 51: 	119 
    -- CP-element group 51: 	156 
    -- CP-element group 51: 	157 
    -- CP-element group 51: 	167 
    -- CP-element group 51: 	169 
    -- CP-element group 51: 	186 
    -- CP-element group 51: 	214 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/loop_body_start
      -- CP-element group 51: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/$entry
      -- 
    -- Element group convTransposeC_CP_5701_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	213 
    -- CP-element group 52: 	214 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	47 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/condition_evaluated
      -- 
    condition_evaluated_6025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(52), ack => do_while_stmt_2389_branch_req_0); -- 
    convTransposeC_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(56) & convTransposeC_CP_5701_elements(213) & convTransposeC_CP_5701_elements(214);
      gj_convTransposeC_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	57 
    -- CP-element group 53: 	76 
    -- CP-element group 53: 	97 
    -- CP-element group 53: 	118 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53: 	99 
    -- CP-element group 53: 	120 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/aggregated_phi_sample_req
      -- CP-element group 53: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_sample_start__ps
      -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(57) & convTransposeC_CP_5701_elements(76) & convTransposeC_CP_5701_elements(97) & convTransposeC_CP_5701_elements(118) & convTransposeC_CP_5701_elements(56);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	59 
    -- CP-element group 54: 	79 
    -- CP-element group 54: 	100 
    -- CP-element group 54: 	121 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	183 
    -- CP-element group 54: 	187 
    -- CP-element group 54: 	191 
    -- CP-element group 54: 	195 
    -- CP-element group 54: 	199 
    -- CP-element group 54: 	203 
    -- CP-element group 54: 	207 
    -- CP-element group 54: 	215 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: 	76 
    -- CP-element group 54: 	97 
    -- CP-element group 54: 	118 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/aggregated_phi_sample_ack
      -- CP-element group 54: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_sample_completed_
      -- 
    convTransposeC_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(59) & convTransposeC_CP_5701_elements(79) & convTransposeC_CP_5701_elements(100) & convTransposeC_CP_5701_elements(121);
      gj_convTransposeC_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	77 
    -- CP-element group 55: 	98 
    -- CP-element group 55: 	119 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	80 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	122 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/aggregated_phi_update_req
      -- CP-element group 55: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_update_start__ps
      -- 
    convTransposeC_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(58) & convTransposeC_CP_5701_elements(77) & convTransposeC_CP_5701_elements(98) & convTransposeC_CP_5701_elements(119);
      gj_convTransposeC_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	81 
    -- CP-element group 56: 	102 
    -- CP-element group 56: 	123 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/aggregated_phi_update_ack
      -- 
    convTransposeC_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(60) & convTransposeC_CP_5701_elements(81) & convTransposeC_CP_5701_elements(102) & convTransposeC_CP_5701_elements(123);
      gj_convTransposeC_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	53 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_sample_start_
      -- 
    convTransposeC_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(54);
      gj_convTransposeC_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	153 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	55 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_update_start_
      -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(60) & convTransposeC_CP_5701_elements(153);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	54 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_sample_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: 	151 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_update_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	49 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_loopback_trigger
      -- 
    convTransposeC_CP_5701_elements(61) <= convTransposeC_CP_5701_elements(49);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_loopback_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_loopback_sample_req
      -- 
    phi_stmt_2391_loopback_sample_req_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2391_loopback_sample_req_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(62), ack => phi_stmt_2391_req_0); -- 
    -- Element group convTransposeC_CP_5701_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	50 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_entry_trigger
      -- 
    convTransposeC_CP_5701_elements(63) <= convTransposeC_CP_5701_elements(50);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_entry_sample_req_ps
      -- CP-element group 64: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_entry_sample_req
      -- 
    phi_stmt_2391_entry_sample_req_6043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2391_entry_sample_req_6043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(64), ack => phi_stmt_2391_req_1); -- 
    -- Element group convTransposeC_CP_5701_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_phi_mux_ack_ps
      -- CP-element group 65: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2391_phi_mux_ack
      -- 
    phi_stmt_2391_phi_mux_ack_6046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2391_ack_0, ack => convTransposeC_CP_5701_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_sample_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_update_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_sample_start_
      -- 
    rr_6059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(68), ack => type_cast_2394_inst_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(66) & convTransposeC_CP_5701_elements(70);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_update_start_
      -- 
    cr_6064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(69), ack => type_cast_2394_inst_req_1); -- 
    convTransposeC_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(67) & convTransposeC_CP_5701_elements(71);
      gj_convTransposeC_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_sample_completed__ps
      -- 
    ra_6060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2394_inst_ack_0, ack => convTransposeC_CP_5701_elements(70)); -- 
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2394_update_completed__ps
      -- 
    ca_6065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2394_inst_ack_1, ack => convTransposeC_CP_5701_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_sample_start_
      -- 
    -- Element group convTransposeC_CP_5701_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_update_start_
      -- 
    -- Element group convTransposeC_CP_5701_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_update_completed__ps
      -- 
    convTransposeC_CP_5701_elements(74) <= convTransposeC_CP_5701_elements(75);
    -- CP-element group 75:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	74 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_indvar_at_entry_2395_update_completed_
      -- 
    -- Element group convTransposeC_CP_5701_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeC_CP_5701_elements(73), ack => convTransposeC_CP_5701_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	51 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	54 
    -- CP-element group 76: 	185 
    -- CP-element group 76: 	189 
    -- CP-element group 76: 	193 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	53 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_sample_start_
      -- 
    convTransposeC_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(185) & convTransposeC_CP_5701_elements(189) & convTransposeC_CP_5701_elements(193);
      gj_convTransposeC_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	51 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: 	141 
    -- CP-element group 77: 	184 
    -- CP-element group 77: 	192 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	55 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_update_start_
      -- 
    convTransposeC_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(81) & convTransposeC_CP_5701_elements(141) & convTransposeC_CP_5701_elements(184) & convTransposeC_CP_5701_elements(192);
      gj_convTransposeC_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	53 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_sample_start__ps
      -- 
    convTransposeC_CP_5701_elements(78) <= convTransposeC_CP_5701_elements(53);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	54 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_sample_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	55 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_update_start__ps
      -- 
    convTransposeC_CP_5701_elements(80) <= convTransposeC_CP_5701_elements(55);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	56 
    -- CP-element group 81: 	139 
    -- CP-element group 81: 	182 
    -- CP-element group 81: 	190 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_update_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	49 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_loopback_trigger
      -- 
    convTransposeC_CP_5701_elements(82) <= convTransposeC_CP_5701_elements(49);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_loopback_sample_req_ps
      -- 
    phi_stmt_2396_loopback_sample_req_6084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2396_loopback_sample_req_6084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(83), ack => phi_stmt_2396_req_0); -- 
    -- Element group convTransposeC_CP_5701_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	50 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_entry_trigger
      -- 
    convTransposeC_CP_5701_elements(84) <= convTransposeC_CP_5701_elements(50);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_entry_sample_req_ps
      -- CP-element group 85: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_entry_sample_req
      -- 
    phi_stmt_2396_entry_sample_req_6087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2396_entry_sample_req_6087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(85), ack => phi_stmt_2396_req_1); -- 
    -- Element group convTransposeC_CP_5701_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_phi_mux_ack
      -- CP-element group 86: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2396_phi_mux_ack_ps
      -- 
    phi_stmt_2396_phi_mux_ack_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2396_ack_0, ack => convTransposeC_CP_5701_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_sample_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_update_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Sample/$entry
      -- 
    rr_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(89), ack => type_cast_2399_inst_req_0); -- 
    convTransposeC_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(87) & convTransposeC_CP_5701_elements(91);
      gj_convTransposeC_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_update_start_
      -- CP-element group 90: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Update/$entry
      -- 
    cr_6108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(90), ack => type_cast_2399_inst_req_1); -- 
    convTransposeC_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(88) & convTransposeC_CP_5701_elements(92);
      gj_convTransposeC_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Sample/$exit
      -- 
    ra_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_0, ack => convTransposeC_CP_5701_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2399_update_completed_
      -- 
    ca_6109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_1, ack => convTransposeC_CP_5701_elements(92)); -- 
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_sample_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_sample_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_update_start_
      -- CP-element group 94: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_update_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_update_completed__ps
      -- 
    convTransposeC_CP_5701_elements(95) <= convTransposeC_CP_5701_elements(96);
    -- CP-element group 96:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim2x_x1_at_entry_2400_update_completed_
      -- 
    -- Element group convTransposeC_CP_5701_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeC_CP_5701_elements(94), ack => convTransposeC_CP_5701_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	51 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	54 
    -- CP-element group 97: 	197 
    -- CP-element group 97: 	201 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	53 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_sample_start_
      -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(197) & convTransposeC_CP_5701_elements(201);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	51 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: 	145 
    -- CP-element group 98: 	200 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	55 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_update_start_
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(102) & convTransposeC_CP_5701_elements(145) & convTransposeC_CP_5701_elements(200);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	53 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_sample_start__ps
      -- 
    convTransposeC_CP_5701_elements(99) <= convTransposeC_CP_5701_elements(53);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	54 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_sample_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_update_start__ps
      -- 
    convTransposeC_CP_5701_elements(101) <= convTransposeC_CP_5701_elements(55);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	56 
    -- CP-element group 102: 	143 
    -- CP-element group 102: 	198 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_update_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	49 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_loopback_trigger
      -- 
    convTransposeC_CP_5701_elements(103) <= convTransposeC_CP_5701_elements(49);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_loopback_sample_req
      -- 
    phi_stmt_2401_loopback_sample_req_6128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2401_loopback_sample_req_6128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(104), ack => phi_stmt_2401_req_0); -- 
    -- Element group convTransposeC_CP_5701_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	50 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_entry_trigger
      -- 
    convTransposeC_CP_5701_elements(105) <= convTransposeC_CP_5701_elements(50);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_entry_sample_req
      -- 
    phi_stmt_2401_entry_sample_req_6131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2401_entry_sample_req_6131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(106), ack => phi_stmt_2401_req_1); -- 
    -- Element group convTransposeC_CP_5701_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2401_phi_mux_ack_ps
      -- 
    phi_stmt_2401_phi_mux_ack_6134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2401_ack_0, ack => convTransposeC_CP_5701_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_sample_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_update_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Sample/$entry
      -- 
    rr_6147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(110), ack => type_cast_2404_inst_req_0); -- 
    convTransposeC_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(108) & convTransposeC_CP_5701_elements(112);
      gj_convTransposeC_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_update_start_
      -- 
    cr_6152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(111), ack => type_cast_2404_inst_req_1); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(109) & convTransposeC_CP_5701_elements(113);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Sample/$exit
      -- 
    ra_6148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_0, ack => convTransposeC_CP_5701_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2404_update_completed_
      -- 
    ca_6153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2404_inst_ack_1, ack => convTransposeC_CP_5701_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_sample_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_update_start_
      -- 
    -- Element group convTransposeC_CP_5701_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_update_completed__ps
      -- 
    convTransposeC_CP_5701_elements(116) <= convTransposeC_CP_5701_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim1x_x1_at_entry_2405_update_completed_
      -- 
    -- Element group convTransposeC_CP_5701_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convTransposeC_CP_5701_elements(115), ack => convTransposeC_CP_5701_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	51 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	54 
    -- CP-element group 118: 	205 
    -- CP-element group 118: 	209 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	53 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_sample_start_
      -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(205) & convTransposeC_CP_5701_elements(209);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	51 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	149 
    -- CP-element group 119: 	208 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	55 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_update_start_
      -- 
    convTransposeC_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(123) & convTransposeC_CP_5701_elements(149) & convTransposeC_CP_5701_elements(208);
      gj_convTransposeC_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	53 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_sample_start__ps
      -- 
    convTransposeC_CP_5701_elements(120) <= convTransposeC_CP_5701_elements(53);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	54 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_sample_completed__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	55 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_update_start__ps
      -- 
    convTransposeC_CP_5701_elements(122) <= convTransposeC_CP_5701_elements(55);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	56 
    -- CP-element group 123: 	147 
    -- CP-element group 123: 	206 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	119 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_update_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_update_completed_
      -- 
    -- Element group convTransposeC_CP_5701_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	49 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_loopback_trigger
      -- 
    convTransposeC_CP_5701_elements(124) <= convTransposeC_CP_5701_elements(49);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_loopback_sample_req
      -- CP-element group 125: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_loopback_sample_req_ps
      -- 
    phi_stmt_2406_loopback_sample_req_6172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2406_loopback_sample_req_6172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(125), ack => phi_stmt_2406_req_0); -- 
    -- Element group convTransposeC_CP_5701_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	50 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_entry_trigger
      -- 
    convTransposeC_CP_5701_elements(126) <= convTransposeC_CP_5701_elements(50);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_entry_sample_req_ps
      -- 
    phi_stmt_2406_entry_sample_req_6175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2406_entry_sample_req_6175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(127), ack => phi_stmt_2406_req_1); -- 
    -- Element group convTransposeC_CP_5701_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/phi_stmt_2406_phi_mux_ack_ps
      -- 
    phi_stmt_2406_phi_mux_ack_6178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2406_ack_0, ack => convTransposeC_CP_5701_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_sample_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_update_start__ps
      -- 
    -- Element group convTransposeC_CP_5701_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_sample_start_
      -- 
    rr_6191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(131), ack => type_cast_2409_inst_req_0); -- 
    convTransposeC_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(129) & convTransposeC_CP_5701_elements(133);
      gj_convTransposeC_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_update_start_
      -- CP-element group 132: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Update/cr
      -- 
    cr_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(132), ack => type_cast_2409_inst_req_1); -- 
    convTransposeC_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(130) & convTransposeC_CP_5701_elements(134);
      gj_convTransposeC_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_sample_completed_
      -- 
    ra_6192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_0, ack => convTransposeC_CP_5701_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2409_Update/ca
      -- 
    ca_6197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_1, ack => convTransposeC_CP_5701_elements(134)); -- 
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Sample/req
      -- CP-element group 135: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_sample_start__ps
      -- 
    req_6209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(135), ack => input_dim0x_x1_at_entry_2384_2410_buf_req_0); -- 
    -- Element group convTransposeC_CP_5701_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_update_start_
      -- CP-element group 136: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_update_start__ps
      -- CP-element group 136: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Update/req
      -- 
    req_6214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(136), ack => input_dim0x_x1_at_entry_2384_2410_buf_req_1); -- 
    -- Element group convTransposeC_CP_5701_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_sample_completed__ps
      -- 
    ack_6210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_dim0x_x1_at_entry_2384_2410_buf_ack_0, ack => convTransposeC_CP_5701_elements(137)); -- 
    -- CP-element group 138:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Update/ack
      -- CP-element group 138: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/R_input_dim0x_x1_at_entry_2410_update_completed__ps
      -- 
    ack_6215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_dim0x_x1_at_entry_2384_2410_buf_ack_1, ack => convTransposeC_CP_5701_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	81 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Sample/$entry
      -- 
    rr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(139), ack => type_cast_2439_inst_req_0); -- 
    convTransposeC_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(81) & convTransposeC_CP_5701_elements(141);
      gj_convTransposeC_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: 	170 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_update_start_
      -- CP-element group 140: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Update/cr
      -- 
    cr_6229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(140), ack => type_cast_2439_inst_req_1); -- 
    convTransposeC_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(142) & convTransposeC_CP_5701_elements(170);
      gj_convTransposeC_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	77 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_sample_completed_
      -- 
    ra_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2439_inst_ack_0, ack => convTransposeC_CP_5701_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	168 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2439_update_completed_
      -- 
    ca_6230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2439_inst_ack_1, ack => convTransposeC_CP_5701_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	102 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_sample_start_
      -- 
    rr_6238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(143), ack => type_cast_2443_inst_req_0); -- 
    convTransposeC_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(102) & convTransposeC_CP_5701_elements(145);
      gj_convTransposeC_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: 	170 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_update_start_
      -- CP-element group 144: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Update/cr
      -- 
    cr_6243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(144), ack => type_cast_2443_inst_req_1); -- 
    convTransposeC_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(146) & convTransposeC_CP_5701_elements(170);
      gj_convTransposeC_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	98 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Sample/ra
      -- 
    ra_6239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2443_inst_ack_0, ack => convTransposeC_CP_5701_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	168 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2443_Update/$exit
      -- 
    ca_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2443_inst_ack_1, ack => convTransposeC_CP_5701_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	123 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_sample_start_
      -- 
    rr_6252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(147), ack => type_cast_2447_inst_req_0); -- 
    convTransposeC_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(123) & convTransposeC_CP_5701_elements(149);
      gj_convTransposeC_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: 	170 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Update/cr
      -- CP-element group 148: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_update_start_
      -- 
    cr_6257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(148), ack => type_cast_2447_inst_req_1); -- 
    convTransposeC_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(150) & convTransposeC_CP_5701_elements(170);
      gj_convTransposeC_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	119 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_sample_completed_
      -- 
    ra_6253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2447_inst_ack_0, ack => convTransposeC_CP_5701_elements(149)); -- 
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	168 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2447_Update/ca
      -- 
    ca_6258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2447_inst_ack_1, ack => convTransposeC_CP_5701_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	60 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Sample/rr
      -- 
    rr_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(151), ack => type_cast_2471_inst_req_0); -- 
    convTransposeC_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(60) & convTransposeC_CP_5701_elements(153);
      gj_convTransposeC_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: 	158 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_update_start_
      -- CP-element group 152: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Update/cr
      -- 
    cr_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(152), ack => type_cast_2471_inst_req_1); -- 
    convTransposeC_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(154) & convTransposeC_CP_5701_elements(158);
      gj_convTransposeC_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	58 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Sample/ra
      -- 
    ra_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2471_inst_ack_0, ack => convTransposeC_CP_5701_elements(153)); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	158 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (16) 
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2471_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_resized_1
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_scaled_1
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_computed_1
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_resize_1/$entry
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_resize_1/$exit
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_resize_1/index_resize_req
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_resize_1/index_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_scale_1/$entry
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_scale_1/$exit
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_scale_1/scale_rename_req
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_index_scale_1/scale_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Sample/req
      -- 
    ca_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2471_inst_ack_1, ack => convTransposeC_CP_5701_elements(154)); -- 
    req_6297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(154), ack => array_obj_ref_2477_index_offset_req_0); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	160 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	160 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_request/$entry
      -- CP-element group 155: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_request/req
      -- 
    req_6312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(155), ack => addr_of_2478_final_reg_req_0); -- 
    convTransposeC_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(159) & convTransposeC_CP_5701_elements(160);
      gj_convTransposeC_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	51 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	164 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_update_start_
      -- CP-element group 156: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_complete/req
      -- 
    req_6317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(156), ack => addr_of_2478_final_reg_req_1); -- 
    convTransposeC_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(161) & convTransposeC_CP_5701_elements(164);
      gj_convTransposeC_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	51 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_update_start
      -- CP-element group 157: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Update/req
      -- 
    req_6302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(157), ack => array_obj_ref_2477_index_offset_req_1); -- 
    convTransposeC_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(159) & convTransposeC_CP_5701_elements(160);
      gj_convTransposeC_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	215 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	152 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_sample_complete
      -- CP-element group 158: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Sample/ack
      -- 
    ack_6298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2477_index_offset_ack_0, ack => convTransposeC_CP_5701_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (8) 
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_root_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_offset_calculated
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_final_index_sum_regn_Update/ack
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_base_plus_offset/$entry
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_base_plus_offset/$exit
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_base_plus_offset/sum_rename_req
      -- CP-element group 159: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2477_base_plus_offset/sum_rename_ack
      -- 
    ack_6303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2477_index_offset_ack_1, ack => convTransposeC_CP_5701_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_request/$exit
      -- CP-element group 160: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_request/ack
      -- 
    ack_6313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2478_final_reg_ack_0, ack => convTransposeC_CP_5701_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (19) 
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_complete/$exit
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2478_complete/ack
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_word_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_root_address_calculated
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_address_resized
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_addr_resize/$entry
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_addr_resize/$exit
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_addr_resize/base_resize_req
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_addr_resize/base_resize_ack
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_plus_offset/$entry
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_plus_offset/$exit
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_plus_offset/sum_rename_req
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_base_plus_offset/sum_rename_ack
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_word_addrgen/$entry
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_word_addrgen/$exit
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_word_addrgen/root_register_req
      -- CP-element group 161: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_word_addrgen/root_register_ack
      -- 
    ack_6318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2478_final_reg_ack_1, ack => convTransposeC_CP_5701_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/word_access_start/word_0/rr
      -- 
    rr_6351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(162), ack => ptr_deref_2482_load_0_req_0); -- 
    convTransposeC_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(161) & convTransposeC_CP_5701_elements(164);
      gj_convTransposeC_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: 	180 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_update_start_
      -- CP-element group 163: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/word_access_complete/word_0/cr
      -- 
    cr_6362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(163), ack => ptr_deref_2482_load_0_req_1); -- 
    convTransposeC_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(165) & convTransposeC_CP_5701_elements(180);
      gj_convTransposeC_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/word_access_start/$exit
      -- CP-element group 164: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/word_access_start/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Sample/word_access_start/word_0/ra
      -- 
    ra_6352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2482_load_0_ack_0, ack => convTransposeC_CP_5701_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	178 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (9) 
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/word_access_complete/$exit
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/word_access_complete/word_0/$exit
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/word_access_complete/word_0/ca
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/ptr_deref_2482_Merge/$entry
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/ptr_deref_2482_Merge/$exit
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/ptr_deref_2482_Merge/merge_req
      -- CP-element group 165: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2482_Update/ptr_deref_2482_Merge/merge_ack
      -- 
    ca_6363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2482_load_0_ack_1, ack => convTransposeC_CP_5701_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	171 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	172 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	172 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_request/$entry
      -- CP-element group 166: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_request/req
      -- 
    req_6408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(166), ack => addr_of_2501_final_reg_req_0); -- 
    convTransposeC_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(171) & convTransposeC_CP_5701_elements(172);
      gj_convTransposeC_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	51 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	173 
    -- CP-element group 167: 	176 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	173 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_complete/req
      -- 
    req_6413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(167), ack => addr_of_2501_final_reg_req_1); -- 
    convTransposeC_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(173) & convTransposeC_CP_5701_elements(176);
      gj_convTransposeC_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	142 
    -- CP-element group 168: 	146 
    -- CP-element group 168: 	150 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (13) 
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_resized_1
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_scaled_1
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_computed_1
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_resize_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_resize_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_resize_1/index_resize_req
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_resize_1/index_resize_ack
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_scale_1/$entry
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_scale_1/$exit
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_scale_1/scale_rename_req
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_index_scale_1/scale_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Sample/req
      -- 
    req_6393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(168), ack => array_obj_ref_2500_index_offset_req_0); -- 
    convTransposeC_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(142) & convTransposeC_CP_5701_elements(146) & convTransposeC_CP_5701_elements(150);
      gj_convTransposeC_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	51 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_update_start
      -- CP-element group 169: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Update/req
      -- 
    req_6398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(169), ack => array_obj_ref_2500_index_offset_req_1); -- 
    convTransposeC_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(171) & convTransposeC_CP_5701_elements(172);
      gj_convTransposeC_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	215 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	140 
    -- CP-element group 170: 	144 
    -- CP-element group 170: 	148 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_sample_complete
      -- CP-element group 170: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Sample/ack
      -- 
    ack_6394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2500_index_offset_ack_0, ack => convTransposeC_CP_5701_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	166 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (8) 
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/array_obj_ref_2500_base_plus_offset/sum_rename_ack
      -- 
    ack_6399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2500_index_offset_ack_1, ack => convTransposeC_CP_5701_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_request/$exit
      -- CP-element group 172: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_request/ack
      -- 
    ack_6409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2501_final_reg_ack_0, ack => convTransposeC_CP_5701_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	167 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	167 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/addr_of_2501_complete/ack
      -- 
    ack_6414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2501_final_reg_ack_1, ack => convTransposeC_CP_5701_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Sample/req
      -- 
    req_6422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(174), ack => W_arrayidx86_2473_delayed_6_0_2503_inst_req_0); -- 
    convTransposeC_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(173) & convTransposeC_CP_5701_elements(176);
      gj_convTransposeC_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: 	180 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_update_start_
      -- CP-element group 175: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Update/req
      -- 
    req_6427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(175), ack => W_arrayidx86_2473_delayed_6_0_2503_inst_req_1); -- 
    convTransposeC_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(177) & convTransposeC_CP_5701_elements(180);
      gj_convTransposeC_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	167 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Sample/ack
      -- 
    ack_6423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx86_2473_delayed_6_0_2503_inst_ack_0, ack => convTransposeC_CP_5701_elements(176)); -- 
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (19) 
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2505_Update/ack
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_word_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_root_address_calculated
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_address_resized
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_addr_resize/$entry
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_addr_resize/$exit
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_addr_resize/base_resize_req
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_addr_resize/base_resize_ack
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_plus_offset/$entry
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_plus_offset/$exit
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_plus_offset/sum_rename_req
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_base_plus_offset/sum_rename_ack
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_word_addrgen/$entry
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_word_addrgen/$exit
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_word_addrgen/root_register_req
      -- CP-element group 177: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_word_addrgen/root_register_ack
      -- 
    ack_6428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx86_2473_delayed_6_0_2503_inst_ack_1, ack => convTransposeC_CP_5701_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	165 
    -- CP-element group 178: 	177 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/ptr_deref_2507_Split/$entry
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/ptr_deref_2507_Split/$exit
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/ptr_deref_2507_Split/split_req
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/ptr_deref_2507_Split/split_ack
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/word_access_start/$entry
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/word_access_start/word_0/$entry
      -- CP-element group 178: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/word_access_start/word_0/rr
      -- 
    rr_6466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(178), ack => ptr_deref_2507_store_0_req_0); -- 
    convTransposeC_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(165) & convTransposeC_CP_5701_elements(177) & convTransposeC_CP_5701_elements(180);
      gj_convTransposeC_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (5) 
      -- CP-element group 179: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_update_start_
      -- CP-element group 179: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/word_access_complete/$entry
      -- CP-element group 179: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/word_access_complete/word_0/$entry
      -- CP-element group 179: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/word_access_complete/word_0/cr
      -- 
    cr_6477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(179), ack => ptr_deref_2507_store_0_req_1); -- 
    convTransposeC_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeC_CP_5701_elements(181);
      gj_convTransposeC_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	163 
    -- CP-element group 180: 	175 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/word_access_start/$exit
      -- CP-element group 180: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/word_access_start/word_0/$exit
      -- CP-element group 180: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Sample/word_access_start/word_0/ra
      -- 
    ra_6467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2507_store_0_ack_0, ack => convTransposeC_CP_5701_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	215 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/word_access_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/word_access_complete/word_0/$exit
      -- CP-element group 181: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/ptr_deref_2507_Update/word_access_complete/word_0/ca
      -- 
    ca_6478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2507_store_0_ack_1, ack => convTransposeC_CP_5701_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	81 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Sample/rr
      -- 
    rr_6486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(182), ack => type_cast_2512_inst_req_0); -- 
    convTransposeC_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(81) & convTransposeC_CP_5701_elements(184);
      gj_convTransposeC_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	54 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: 	196 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_update_start_
      -- CP-element group 183: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Update/cr
      -- 
    cr_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(183), ack => type_cast_2512_inst_req_1); -- 
    convTransposeC_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(185) & convTransposeC_CP_5701_elements(196);
      gj_convTransposeC_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	77 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Sample/ra
      -- 
    ra_6487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_0, ack => convTransposeC_CP_5701_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	194 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	76 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2512_Update/ca
      -- 
    ca_6492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_1, ack => convTransposeC_CP_5701_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	51 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Sample/rr
      -- 
    rr_6500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(186), ack => type_cast_2516_inst_req_0); -- 
    convTransposeC_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(51) & convTransposeC_CP_5701_elements(188);
      gj_convTransposeC_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	54 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	189 
    -- CP-element group 187: 	196 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_update_start_
      -- CP-element group 187: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Update/cr
      -- 
    cr_6505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(187), ack => type_cast_2516_inst_req_1); -- 
    convTransposeC_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(189) & convTransposeC_CP_5701_elements(196);
      gj_convTransposeC_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Sample/ra
      -- 
    ra_6501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2516_inst_ack_0, ack => convTransposeC_CP_5701_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	194 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	76 
    -- CP-element group 189: 	187 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2516_Update/ca
      -- 
    ca_6506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2516_inst_ack_1, ack => convTransposeC_CP_5701_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	81 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Sample/req
      -- 
    req_6514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(190), ack => W_add101_2496_delayed_1_0_2530_inst_req_0); -- 
    convTransposeC_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(81) & convTransposeC_CP_5701_elements(192);
      gj_convTransposeC_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	54 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_update_start_
      -- CP-element group 191: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Update/req
      -- 
    req_6519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(191), ack => W_add101_2496_delayed_1_0_2530_inst_req_1); -- 
    convTransposeC_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(193);
      gj_convTransposeC_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	77 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Sample/ack
      -- 
    ack_6515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add101_2496_delayed_1_0_2530_inst_ack_0, ack => convTransposeC_CP_5701_elements(192)); -- 
    -- CP-element group 193:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	215 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	76 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2532_Update/ack
      -- 
    ack_6520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add101_2496_delayed_1_0_2530_inst_ack_1, ack => convTransposeC_CP_5701_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	185 
    -- CP-element group 194: 	189 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Sample/rr
      -- 
    rr_6528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(194), ack => type_cast_2542_inst_req_0); -- 
    convTransposeC_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(185) & convTransposeC_CP_5701_elements(189) & convTransposeC_CP_5701_elements(196);
      gj_convTransposeC_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	54 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: 	204 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_update_start_
      -- CP-element group 195: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Update/cr
      -- 
    cr_6533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(195), ack => type_cast_2542_inst_req_1); -- 
    convTransposeC_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(197) & convTransposeC_CP_5701_elements(204);
      gj_convTransposeC_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	183 
    -- CP-element group 196: 	187 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Sample/ra
      -- 
    ra_6529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2542_inst_ack_0, ack => convTransposeC_CP_5701_elements(196)); -- 
    -- CP-element group 197:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	202 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	97 
    -- CP-element group 197: 	195 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2542_Update/ca
      -- 
    ca_6534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2542_inst_ack_1, ack => convTransposeC_CP_5701_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	102 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Sample/req
      -- 
    req_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(198), ack => W_input_dim1x_x1_2513_delayed_2_0_2550_inst_req_0); -- 
    convTransposeC_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(102) & convTransposeC_CP_5701_elements(200);
      gj_convTransposeC_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	54 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	201 
    -- CP-element group 199: 	204 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_update_start_
      -- CP-element group 199: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Update/req
      -- 
    req_6547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(199), ack => W_input_dim1x_x1_2513_delayed_2_0_2550_inst_req_1); -- 
    convTransposeC_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(201) & convTransposeC_CP_5701_elements(204);
      gj_convTransposeC_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	98 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Sample/ack
      -- 
    ack_6543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_2513_delayed_2_0_2550_inst_ack_0, ack => convTransposeC_CP_5701_elements(200)); -- 
    -- CP-element group 201:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	97 
    -- CP-element group 201: 	199 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2552_Update/ack
      -- 
    ack_6548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_2513_delayed_2_0_2550_inst_ack_1, ack => convTransposeC_CP_5701_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	197 
    -- CP-element group 202: 	201 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Sample/rr
      -- 
    rr_6556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(202), ack => type_cast_2565_inst_req_0); -- 
    convTransposeC_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(197) & convTransposeC_CP_5701_elements(201) & convTransposeC_CP_5701_elements(204);
      gj_convTransposeC_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	54 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: 	212 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_update_start_
      -- CP-element group 203: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Update/cr
      -- 
    cr_6561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(203), ack => type_cast_2565_inst_req_1); -- 
    convTransposeC_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(205) & convTransposeC_CP_5701_elements(212);
      gj_convTransposeC_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	195 
    -- CP-element group 204: 	199 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Sample/ra
      -- 
    ra_6557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_0, ack => convTransposeC_CP_5701_elements(204)); -- 
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	210 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	118 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2565_Update/ca
      -- 
    ca_6562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2565_inst_ack_1, ack => convTransposeC_CP_5701_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	123 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Sample/req
      -- 
    req_6570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(206), ack => W_input_dim0x_x1_2527_delayed_3_0_2567_inst_req_0); -- 
    convTransposeC_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(123) & convTransposeC_CP_5701_elements(208);
      gj_convTransposeC_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	54 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: 	212 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_update_start_
      -- CP-element group 207: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Update/req
      -- 
    req_6575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(207), ack => W_input_dim0x_x1_2527_delayed_3_0_2567_inst_req_1); -- 
    convTransposeC_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(209) & convTransposeC_CP_5701_elements(212);
      gj_convTransposeC_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	119 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Sample/ack
      -- 
    ack_6571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_2527_delayed_3_0_2567_inst_ack_0, ack => convTransposeC_CP_5701_elements(208)); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	118 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/assign_stmt_2569_Update/ack
      -- 
    ack_6576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_2527_delayed_3_0_2567_inst_ack_1, ack => convTransposeC_CP_5701_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	205 
    -- CP-element group 210: 	209 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Sample/rr
      -- 
    rr_6584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(210), ack => type_cast_2584_inst_req_0); -- 
    convTransposeC_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(205) & convTransposeC_CP_5701_elements(209) & convTransposeC_CP_5701_elements(212);
      gj_convTransposeC_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_update_start_
      -- CP-element group 211: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Update/cr
      -- 
    cr_6589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(211), ack => type_cast_2584_inst_req_1); -- 
    convTransposeC_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeC_CP_5701_elements(213);
      gj_convTransposeC_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	203 
    -- CP-element group 212: 	207 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Sample/ra
      -- 
    ra_6585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2584_inst_ack_0, ack => convTransposeC_CP_5701_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	52 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/type_cast_2584_Update/ca
      -- 
    ca_6590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2584_inst_ack_1, ack => convTransposeC_CP_5701_elements(213)); -- 
    -- CP-element group 214:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	51 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	52 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convTransposeC_CP_5701_elements(214) is a control-delay.
    cp_element_214_delay: control_delay_element  generic map(name => " 214_delay", delay_value => 1)  port map(req => convTransposeC_CP_5701_elements(51), ack => convTransposeC_CP_5701_elements(214), clk => clk, reset =>reset);
    -- CP-element group 215:  join  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	54 
    -- CP-element group 215: 	158 
    -- CP-element group 215: 	170 
    -- CP-element group 215: 	181 
    -- CP-element group 215: 	193 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	48 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_2236/do_while_stmt_2389/do_while_stmt_2389_loop_body/$exit
      -- 
    convTransposeC_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(54) & convTransposeC_CP_5701_elements(158) & convTransposeC_CP_5701_elements(170) & convTransposeC_CP_5701_elements(181) & convTransposeC_CP_5701_elements(193);
      gj_convTransposeC_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_exit/$exit
      -- CP-element group 216: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_exit/ack
      -- 
    ack_6595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2389_branch_ack_0, ack => convTransposeC_CP_5701_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	47 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_taken/$exit
      -- CP-element group 217: 	 branch_block_stmt_2236/do_while_stmt_2389/loop_taken/ack
      -- 
    ack_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2389_branch_ack_1, ack => convTransposeC_CP_5701_elements(217)); -- 
    -- CP-element group 218:  transition  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	1 
    -- CP-element group 218:  members (1) 
      -- CP-element group 218: 	 branch_block_stmt_2236/do_while_stmt_2389/$exit
      -- 
    convTransposeC_CP_5701_elements(218) <= convTransposeC_CP_5701_elements(45);
    -- CP-element group 219:  merge  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	1 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (15) 
      -- CP-element group 219: 	 branch_block_stmt_2236/merge_stmt_2607__exit__
      -- CP-element group 219: 	 branch_block_stmt_2236/assign_stmt_2612__entry__
      -- CP-element group 219: 	 branch_block_stmt_2236/if_stmt_2603_if_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_2236/if_stmt_2603_if_link/if_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_2236/whilex_xbody_whilex_xend
      -- CP-element group 219: 	 branch_block_stmt_2236/assign_stmt_2612/$entry
      -- CP-element group 219: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Sample/req
      -- CP-element group 219: 	 branch_block_stmt_2236/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_2236/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_2236/merge_stmt_2607_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_2236/merge_stmt_2607_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_2236/merge_stmt_2607_PhiAck/$exit
      -- CP-element group 219: 	 branch_block_stmt_2236/merge_stmt_2607_PhiAck/dummy
      -- 
    if_choice_transition_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2603_branch_ack_1, ack => convTransposeC_CP_5701_elements(219)); -- 
    req_6629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(219), ack => WPIPE_Block2_done_2609_inst_req_0); -- 
    -- CP-element group 220:  merge  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	1 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_2236/if_stmt_2603__exit__
      -- CP-element group 220: 	 branch_block_stmt_2236/merge_stmt_2607__entry__
      -- CP-element group 220: 	 branch_block_stmt_2236/if_stmt_2603_else_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_2236/if_stmt_2603_else_link/else_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_2236/merge_stmt_2607_dead_link/$entry
      -- 
    else_choice_transition_6617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2603_branch_ack_0, ack => convTransposeC_CP_5701_elements(220)); -- 
    -- CP-element group 221:  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_update_start_
      -- CP-element group 221: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Sample/ack
      -- CP-element group 221: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Update/req
      -- 
    ack_6630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2609_inst_ack_0, ack => convTransposeC_CP_5701_elements(221)); -- 
    req_6634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(221), ack => WPIPE_Block2_done_2609_inst_req_1); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (16) 
      -- CP-element group 222: 	 $exit
      -- CP-element group 222: 	 branch_block_stmt_2236/$exit
      -- CP-element group 222: 	 branch_block_stmt_2236/branch_block_stmt_2236__exit__
      -- CP-element group 222: 	 branch_block_stmt_2236/assign_stmt_2612__exit__
      -- CP-element group 222: 	 branch_block_stmt_2236/return__
      -- CP-element group 222: 	 branch_block_stmt_2236/merge_stmt_2614__exit__
      -- CP-element group 222: 	 branch_block_stmt_2236/assign_stmt_2612/$exit
      -- CP-element group 222: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_2236/assign_stmt_2612/WPIPE_Block2_done_2609_Update/ack
      -- CP-element group 222: 	 branch_block_stmt_2236/return___PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_2236/return___PhiReq/$exit
      -- CP-element group 222: 	 branch_block_stmt_2236/merge_stmt_2614_PhiReqMerge
      -- CP-element group 222: 	 branch_block_stmt_2236/merge_stmt_2614_PhiAck/$entry
      -- CP-element group 222: 	 branch_block_stmt_2236/merge_stmt_2614_PhiAck/$exit
      -- CP-element group 222: 	 branch_block_stmt_2236/merge_stmt_2614_PhiAck/dummy
      -- 
    ack_6635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2609_inst_ack_1, ack => convTransposeC_CP_5701_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	43 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Sample/ra
      -- 
    ra_6655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2387_inst_ack_0, ack => convTransposeC_CP_5701_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	43 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/Update/ca
      -- 
    ca_6660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2387_inst_ack_1, ack => convTransposeC_CP_5701_elements(224)); -- 
    -- CP-element group 225:  join  transition  place  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (8) 
      -- CP-element group 225: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/$exit
      -- CP-element group 225: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/$exit
      -- CP-element group 225: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/$exit
      -- CP-element group 225: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/$exit
      -- CP-element group 225: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_sources/type_cast_2387/SplitProtocol/$exit
      -- CP-element group 225: 	 branch_block_stmt_2236/entry_whilex_xbody_PhiReq/phi_stmt_2384/phi_stmt_2384_req
      -- CP-element group 225: 	 branch_block_stmt_2236/merge_stmt_2368_PhiReqMerge
      -- CP-element group 225: 	 branch_block_stmt_2236/merge_stmt_2368_PhiAck/$entry
      -- 
    phi_stmt_2384_req_6661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2384_req_6661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5701_elements(225), ack => phi_stmt_2384_req_0); -- 
    convTransposeC_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5701_elements(223) & convTransposeC_CP_5701_elements(224);
      gj_convTransposeC_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5701_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  transition  place  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	44 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_2236/merge_stmt_2368__exit__
      -- CP-element group 226: 	 branch_block_stmt_2236/do_while_stmt_2389__entry__
      -- CP-element group 226: 	 branch_block_stmt_2236/merge_stmt_2368_PhiAck/$exit
      -- CP-element group 226: 	 branch_block_stmt_2236/merge_stmt_2368_PhiAck/phi_stmt_2384_ack
      -- 
    phi_stmt_2384_ack_6666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2384_ack_0, ack => convTransposeC_CP_5701_elements(226)); -- 
    convTransposeC_do_while_stmt_2389_terminator_6600: loop_terminator -- 
      generic map (name => " convTransposeC_do_while_stmt_2389_terminator_6600", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convTransposeC_CP_5701_elements(48),loop_continue => convTransposeC_CP_5701_elements(217),loop_terminate => convTransposeC_CP_5701_elements(216),loop_back => convTransposeC_CP_5701_elements(46),loop_exit => convTransposeC_CP_5701_elements(45),clk => clk, reset => reset); -- 
    phi_stmt_2391_phi_seq_6074_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeC_CP_5701_elements(61);
      convTransposeC_CP_5701_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeC_CP_5701_elements(70);
      convTransposeC_CP_5701_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeC_CP_5701_elements(71);
      convTransposeC_CP_5701_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeC_CP_5701_elements(63);
      convTransposeC_CP_5701_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeC_CP_5701_elements(72);
      convTransposeC_CP_5701_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeC_CP_5701_elements(74);
      convTransposeC_CP_5701_elements(64) <= phi_mux_reqs(1);
      phi_stmt_2391_phi_seq_6074 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2391_phi_seq_6074") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeC_CP_5701_elements(53), 
          phi_sample_ack => convTransposeC_CP_5701_elements(59), 
          phi_update_req => convTransposeC_CP_5701_elements(55), 
          phi_update_ack => convTransposeC_CP_5701_elements(60), 
          phi_mux_ack => convTransposeC_CP_5701_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2396_phi_seq_6118_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeC_CP_5701_elements(82);
      convTransposeC_CP_5701_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeC_CP_5701_elements(91);
      convTransposeC_CP_5701_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeC_CP_5701_elements(92);
      convTransposeC_CP_5701_elements(83) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeC_CP_5701_elements(84);
      convTransposeC_CP_5701_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeC_CP_5701_elements(93);
      convTransposeC_CP_5701_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeC_CP_5701_elements(95);
      convTransposeC_CP_5701_elements(85) <= phi_mux_reqs(1);
      phi_stmt_2396_phi_seq_6118 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2396_phi_seq_6118") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeC_CP_5701_elements(78), 
          phi_sample_ack => convTransposeC_CP_5701_elements(79), 
          phi_update_req => convTransposeC_CP_5701_elements(80), 
          phi_update_ack => convTransposeC_CP_5701_elements(81), 
          phi_mux_ack => convTransposeC_CP_5701_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2401_phi_seq_6162_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeC_CP_5701_elements(103);
      convTransposeC_CP_5701_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeC_CP_5701_elements(112);
      convTransposeC_CP_5701_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeC_CP_5701_elements(113);
      convTransposeC_CP_5701_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeC_CP_5701_elements(105);
      convTransposeC_CP_5701_elements(114)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeC_CP_5701_elements(114);
      convTransposeC_CP_5701_elements(115)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeC_CP_5701_elements(116);
      convTransposeC_CP_5701_elements(106) <= phi_mux_reqs(1);
      phi_stmt_2401_phi_seq_6162 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2401_phi_seq_6162") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeC_CP_5701_elements(99), 
          phi_sample_ack => convTransposeC_CP_5701_elements(100), 
          phi_update_req => convTransposeC_CP_5701_elements(101), 
          phi_update_ack => convTransposeC_CP_5701_elements(102), 
          phi_mux_ack => convTransposeC_CP_5701_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2406_phi_seq_6216_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeC_CP_5701_elements(124);
      convTransposeC_CP_5701_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeC_CP_5701_elements(133);
      convTransposeC_CP_5701_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeC_CP_5701_elements(134);
      convTransposeC_CP_5701_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeC_CP_5701_elements(126);
      convTransposeC_CP_5701_elements(135)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeC_CP_5701_elements(137);
      convTransposeC_CP_5701_elements(136)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeC_CP_5701_elements(138);
      convTransposeC_CP_5701_elements(127) <= phi_mux_reqs(1);
      phi_stmt_2406_phi_seq_6216 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2406_phi_seq_6216") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeC_CP_5701_elements(120), 
          phi_sample_ack => convTransposeC_CP_5701_elements(121), 
          phi_update_req => convTransposeC_CP_5701_elements(122), 
          phi_update_ack => convTransposeC_CP_5701_elements(123), 
          phi_mux_ack => convTransposeC_CP_5701_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6026_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convTransposeC_CP_5701_elements(49);
        preds(1)  <= convTransposeC_CP_5701_elements(50);
        entry_tmerge_6026 : transition_merge -- 
          generic map(name => " entry_tmerge_6026")
          port map (preds => preds, symbol_out => convTransposeC_CP_5701_elements(51));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_2602_wire : std_logic_vector(0 downto 0);
    signal R_idxprom85_2499_resized : std_logic_vector(13 downto 0);
    signal R_idxprom85_2499_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2476_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2476_scaled : std_logic_vector(13 downto 0);
    signal add101_2496_delayed_1_0_2532 : std_logic_vector(15 downto 0);
    signal add101_2529 : std_logic_vector(15 downto 0);
    signal add125_2366 : std_logic_vector(31 downto 0);
    signal add45_2310 : std_logic_vector(15 downto 0);
    signal add58_2321 : std_logic_vector(15 downto 0);
    signal add77_2458 : std_logic_vector(63 downto 0);
    signal add79_2468 : std_logic_vector(63 downto 0);
    signal add_2288 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2416 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2477_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2477_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2500_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2500_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2500_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2500_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2500_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2500_root_address : std_logic_vector(13 downto 0);
    signal arrayidx81_2479 : std_logic_vector(31 downto 0);
    signal arrayidx86_2473_delayed_6_0_2505 : std_logic_vector(31 downto 0);
    signal arrayidx86_2502 : std_logic_vector(31 downto 0);
    signal call11_2257 : std_logic_vector(15 downto 0);
    signal call13_2260 : std_logic_vector(15 downto 0);
    signal call14_2263 : std_logic_vector(15 downto 0);
    signal call15_2266 : std_logic_vector(15 downto 0);
    signal call16_2279 : std_logic_vector(15 downto 0);
    signal call18_2291 : std_logic_vector(15 downto 0);
    signal call1_2242 : std_logic_vector(15 downto 0);
    signal call20_2294 : std_logic_vector(15 downto 0);
    signal call22_2297 : std_logic_vector(15 downto 0);
    signal call3_2245 : std_logic_vector(15 downto 0);
    signal call5_2248 : std_logic_vector(15 downto 0);
    signal call7_2251 : std_logic_vector(15 downto 0);
    signal call9_2254 : std_logic_vector(15 downto 0);
    signal call_2239 : std_logic_vector(15 downto 0);
    signal cmp109_2562 : std_logic_vector(0 downto 0);
    signal cmp126_2590 : std_logic_vector(0 downto 0);
    signal cmp_2523 : std_logic_vector(0 downto 0);
    signal conv116_2585 : std_logic_vector(31 downto 0);
    signal conv119_2349 : std_logic_vector(31 downto 0);
    signal conv17_2283 : std_logic_vector(31 downto 0);
    signal conv65_2440 : std_logic_vector(63 downto 0);
    signal conv68_2330 : std_logic_vector(63 downto 0);
    signal conv70_2444 : std_logic_vector(63 downto 0);
    signal conv73_2334 : std_logic_vector(63 downto 0);
    signal conv75_2448 : std_logic_vector(63 downto 0);
    signal conv95_2513 : std_logic_vector(31 downto 0);
    signal conv97_2345 : std_logic_vector(31 downto 0);
    signal conv_2270 : std_logic_vector(31 downto 0);
    signal iNsTr_18_2543 : std_logic_vector(15 downto 0);
    signal idxprom85_2495 : std_logic_vector(63 downto 0);
    signal idxprom_2472 : std_logic_vector(63 downto 0);
    signal inc113_2566 : std_logic_vector(15 downto 0);
    signal inc113x_xinput_dim0x_x1_2574 : std_logic_vector(15 downto 0);
    signal inc_2549 : std_logic_vector(15 downto 0);
    signal indvar_2391 : std_logic_vector(31 downto 0);
    signal indvar_at_entry_2369 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2596 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1_2406 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_2527_delayed_3_0_2569 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_2384 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_2384_2410_buffered : std_logic_vector(15 downto 0);
    signal input_dim1x_x0_2557 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2401 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2513_delayed_2_0_2552 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_at_entry_2379 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2581 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0_2539 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2396 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_at_entry_2374 : std_logic_vector(15 downto 0);
    signal mul54_2431 : std_logic_vector(15 downto 0);
    signal mul76_2453 : std_logic_vector(63 downto 0);
    signal mul78_2463 : std_logic_vector(63 downto 0);
    signal mul_2421 : std_logic_vector(15 downto 0);
    signal ptr_deref_2482_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2482_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2482_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2482_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2482_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2507_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2507_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2507_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2507_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2507_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2507_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2276 : std_logic_vector(31 downto 0);
    signal shr120140_2355 : std_logic_vector(31 downto 0);
    signal shr124141_2361 : std_logic_vector(31 downto 0);
    signal shr139_2304 : std_logic_vector(15 downto 0);
    signal shr84_2489 : std_logic_vector(63 downto 0);
    signal sub48_2426 : std_logic_vector(15 downto 0);
    signal sub61_2326 : std_logic_vector(15 downto 0);
    signal sub62_2436 : std_logic_vector(15 downto 0);
    signal sub91_2340 : std_logic_vector(15 downto 0);
    signal sub_2315 : std_logic_vector(15 downto 0);
    signal tmp82_2483 : std_logic_vector(63 downto 0);
    signal type_cast_2274_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2302_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2308_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2319_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2338_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2343_wire : std_logic_vector(31 downto 0);
    signal type_cast_2353_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2359_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2387_wire : std_logic_vector(15 downto 0);
    signal type_cast_2394_wire : std_logic_vector(31 downto 0);
    signal type_cast_2399_wire : std_logic_vector(15 downto 0);
    signal type_cast_2404_wire : std_logic_vector(15 downto 0);
    signal type_cast_2409_wire : std_logic_vector(15 downto 0);
    signal type_cast_2485_2485_delayed_2_0_2517 : std_logic_vector(31 downto 0);
    signal type_cast_2487_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2520_wire : std_logic_vector(31 downto 0);
    signal type_cast_2527_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2537_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2547_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2578_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2611_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_whilex_xend_taken_2599 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_2477_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2477_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2477_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2477_resized_base_address <= "00000000000000";
    array_obj_ref_2500_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2500_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2500_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2500_resized_base_address <= "00000000000000";
    indvar_at_entry_2369 <= "00000000000000000000000000000000";
    input_dim1x_x1_at_entry_2379 <= "0000000000000000";
    input_dim2x_x1_at_entry_2374 <= "0000000000000000";
    ptr_deref_2482_word_offset_0 <= "00000000000000";
    ptr_deref_2507_word_offset_0 <= "00000000000000";
    type_cast_2274_wire_constant <= "00000000000000000000000000010000";
    type_cast_2302_wire_constant <= "0000000000000001";
    type_cast_2308_wire_constant <= "1111111111111111";
    type_cast_2319_wire_constant <= "1111111111111111";
    type_cast_2338_wire_constant <= "1111111111111100";
    type_cast_2353_wire_constant <= "00000000000000000000000000000010";
    type_cast_2359_wire_constant <= "00000000000000000000000000000001";
    type_cast_2487_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2493_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2527_wire_constant <= "0000000000000100";
    type_cast_2537_wire_constant <= "0000000000000000";
    type_cast_2547_wire_constant <= "0000000000000001";
    type_cast_2578_wire_constant <= "0000000000000000";
    type_cast_2594_wire_constant <= "00000000000000000000000000000001";
    type_cast_2611_wire_constant <= "0000000000000001";
    phi_stmt_2384: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2387_wire;
      req(0) <= phi_stmt_2384_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2384",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2384_ack_0,
          idata => idata,
          odata => input_dim0x_x1_at_entry_2384,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2384
    phi_stmt_2391: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2394_wire & indvar_at_entry_2369;
      req <= phi_stmt_2391_req_0 & phi_stmt_2391_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2391",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2391_ack_0,
          idata => idata,
          odata => indvar_2391,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2391
    phi_stmt_2396: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2399_wire & input_dim2x_x1_at_entry_2374;
      req <= phi_stmt_2396_req_0 & phi_stmt_2396_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2396",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2396_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2396,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2396
    phi_stmt_2401: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2404_wire & input_dim1x_x1_at_entry_2379;
      req <= phi_stmt_2401_req_0 & phi_stmt_2401_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2401",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2401_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2401,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2401
    phi_stmt_2406: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2409_wire & input_dim0x_x1_at_entry_2384_2410_buffered;
      req <= phi_stmt_2406_req_0 & phi_stmt_2406_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2406",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2406_ack_0,
          idata => idata,
          odata => input_dim0x_x1_2406,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2406
    -- flow-through select operator MUX_2538_inst
    input_dim2x_x0_2539 <= add101_2496_delayed_1_0_2532 when (cmp_2523(0) /=  '0') else type_cast_2537_wire_constant;
    -- flow-through select operator MUX_2580_inst
    input_dim1x_x2_2581 <= type_cast_2578_wire_constant when (cmp109_2562(0) /=  '0') else input_dim1x_x0_2557;
    W_add101_2496_delayed_1_0_2530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add101_2496_delayed_1_0_2530_inst_req_0;
      W_add101_2496_delayed_1_0_2530_inst_ack_0<= wack(0);
      rreq(0) <= W_add101_2496_delayed_1_0_2530_inst_req_1;
      W_add101_2496_delayed_1_0_2530_inst_ack_1<= rack(0);
      W_add101_2496_delayed_1_0_2530_inst : InterlockBuffer generic map ( -- 
        name => "W_add101_2496_delayed_1_0_2530_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add101_2529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add101_2496_delayed_1_0_2532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx86_2473_delayed_6_0_2503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx86_2473_delayed_6_0_2503_inst_req_0;
      W_arrayidx86_2473_delayed_6_0_2503_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx86_2473_delayed_6_0_2503_inst_req_1;
      W_arrayidx86_2473_delayed_6_0_2503_inst_ack_1<= rack(0);
      W_arrayidx86_2473_delayed_6_0_2503_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx86_2473_delayed_6_0_2503_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx86_2502,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_2473_delayed_6_0_2505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim0x_x1_2527_delayed_3_0_2567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim0x_x1_2527_delayed_3_0_2567_inst_req_0;
      W_input_dim0x_x1_2527_delayed_3_0_2567_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim0x_x1_2527_delayed_3_0_2567_inst_req_1;
      W_input_dim0x_x1_2527_delayed_3_0_2567_inst_ack_1<= rack(0);
      W_input_dim0x_x1_2527_delayed_3_0_2567_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim0x_x1_2527_delayed_3_0_2567_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_2406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_2527_delayed_3_0_2569,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim1x_x1_2513_delayed_2_0_2550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim1x_x1_2513_delayed_2_0_2550_inst_req_0;
      W_input_dim1x_x1_2513_delayed_2_0_2550_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim1x_x1_2513_delayed_2_0_2550_inst_req_1;
      W_input_dim1x_x1_2513_delayed_2_0_2550_inst_ack_1<= rack(0);
      W_input_dim1x_x1_2513_delayed_2_0_2550_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim1x_x1_2513_delayed_2_0_2550_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim1x_x1_2513_delayed_2_0_2552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_2597_inst
    process(cmp126_2590) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp126_2590(0 downto 0);
      whilex_xbody_whilex_xend_taken_2599 <= tmp_var; -- 
    end process;
    addr_of_2478_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2478_final_reg_req_0;
      addr_of_2478_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2478_final_reg_req_1;
      addr_of_2478_final_reg_ack_1<= rack(0);
      addr_of_2478_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2478_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2477_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx81_2479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2501_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2501_final_reg_req_0;
      addr_of_2501_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2501_final_reg_req_1;
      addr_of_2501_final_reg_ack_1<= rack(0);
      addr_of_2501_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2501_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2500_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_2502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    input_dim0x_x1_at_entry_2384_2410_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= input_dim0x_x1_at_entry_2384_2410_buf_req_0;
      input_dim0x_x1_at_entry_2384_2410_buf_ack_0<= wack(0);
      rreq(0) <= input_dim0x_x1_at_entry_2384_2410_buf_req_1;
      input_dim0x_x1_at_entry_2384_2410_buf_ack_1<= rack(0);
      input_dim0x_x1_at_entry_2384_2410_buf : InterlockBuffer generic map ( -- 
        name => "input_dim0x_x1_at_entry_2384_2410_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_at_entry_2384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_at_entry_2384_2410_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2269_inst_req_0;
      type_cast_2269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2269_inst_req_1;
      type_cast_2269_inst_ack_1<= rack(0);
      type_cast_2269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2282_inst_req_0;
      type_cast_2282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2282_inst_req_1;
      type_cast_2282_inst_ack_1<= rack(0);
      type_cast_2282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2329_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2329_inst_req_0;
      type_cast_2329_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2329_inst_req_1;
      type_cast_2329_inst_ack_1<= rack(0);
      type_cast_2329_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2329_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2330,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2333_inst_req_0;
      type_cast_2333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2333_inst_req_1;
      type_cast_2333_inst_ack_1<= rack(0);
      type_cast_2333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2344_inst_req_0;
      type_cast_2344_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2344_inst_req_1;
      type_cast_2344_inst_ack_1<= rack(0);
      type_cast_2344_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2344_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2343_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_2345,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2348_inst_req_0;
      type_cast_2348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2348_inst_req_1;
      type_cast_2348_inst_ack_1<= rack(0);
      type_cast_2348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_2349,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2387_inst_req_0;
      type_cast_2387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2387_inst_req_1;
      type_cast_2387_inst_ack_1<= rack(0);
      type_cast_2387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr139_2304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2387_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2394_inst_req_0;
      type_cast_2394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2394_inst_req_1;
      type_cast_2394_inst_ack_1<= rack(0);
      type_cast_2394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2394_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2394_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2399_inst_req_0;
      type_cast_2399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2399_inst_req_1;
      type_cast_2399_inst_ack_1<= rack(0);
      type_cast_2399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2399_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0_2539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2399_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2404_inst_req_0;
      type_cast_2404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2404_inst_req_1;
      type_cast_2404_inst_ack_1<= rack(0);
      type_cast_2404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2404_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2581,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2404_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2409_inst_req_0;
      type_cast_2409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2409_inst_req_1;
      type_cast_2409_inst_ack_1<= rack(0);
      type_cast_2409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2409_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc113x_xinput_dim0x_x1_2574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2409_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2439_inst_req_0;
      type_cast_2439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2439_inst_req_1;
      type_cast_2439_inst_ack_1<= rack(0);
      type_cast_2439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2440,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2443_inst_req_0;
      type_cast_2443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2443_inst_req_1;
      type_cast_2443_inst_ack_1<= rack(0);
      type_cast_2443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2447_inst_req_0;
      type_cast_2447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2447_inst_req_1;
      type_cast_2447_inst_ack_1<= rack(0);
      type_cast_2447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2448,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2471_inst_req_0;
      type_cast_2471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2471_inst_req_1;
      type_cast_2471_inst_ack_1<= rack(0);
      type_cast_2471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_src_0x_x0_2416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2512_inst_req_0;
      type_cast_2512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2512_inst_req_1;
      type_cast_2512_inst_ack_1<= rack(0);
      type_cast_2512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2512_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2516_inst_req_0;
      type_cast_2516_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2516_inst_req_1;
      type_cast_2516_inst_ack_1<= rack(0);
      type_cast_2516_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2516_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv97_2345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2485_2485_delayed_2_0_2517,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2520_inst
    process(conv95_2513) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv95_2513(31 downto 0);
      type_cast_2520_wire <= tmp_var; -- 
    end process;
    type_cast_2542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2542_inst_req_0;
      type_cast_2542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2542_inst_req_1;
      type_cast_2542_inst_ack_1<= rack(0);
      type_cast_2542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2542_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_2523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_18_2543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2565_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2565_inst_req_0;
      type_cast_2565_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2565_inst_req_1;
      type_cast_2565_inst_ack_1<= rack(0);
      type_cast_2565_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2565_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp109_2562,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc113_2566,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2584_inst_req_0;
      type_cast_2584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2584_inst_req_1;
      type_cast_2584_inst_ack_1<= rack(0);
      type_cast_2584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc113x_xinput_dim0x_x1_2574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_2585,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2477_index_1_rename
    process(R_idxprom_2476_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2476_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2476_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2477_index_1_resize
    process(idxprom_2472) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2472;
      ov := iv(13 downto 0);
      R_idxprom_2476_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2477_root_address_inst
    process(array_obj_ref_2477_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2477_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2477_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2500_index_1_rename
    process(R_idxprom85_2499_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom85_2499_resized;
      ov(13 downto 0) := iv;
      R_idxprom85_2499_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2500_index_1_resize
    process(idxprom85_2495) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom85_2495;
      ov := iv(13 downto 0);
      R_idxprom85_2499_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2500_root_address_inst
    process(array_obj_ref_2500_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2500_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2500_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_addr_0
    process(ptr_deref_2482_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2482_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2482_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_base_resize
    process(arrayidx81_2479) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx81_2479;
      ov := iv(13 downto 0);
      ptr_deref_2482_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_gather_scatter
    process(ptr_deref_2482_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2482_data_0;
      ov(63 downto 0) := iv;
      tmp82_2483 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2482_root_address_inst
    process(ptr_deref_2482_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2482_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2482_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2507_addr_0
    process(ptr_deref_2507_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2507_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2507_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2507_base_resize
    process(arrayidx86_2473_delayed_6_0_2505) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx86_2473_delayed_6_0_2505;
      ov := iv(13 downto 0);
      ptr_deref_2507_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2507_gather_scatter
    process(tmp82_2483) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp82_2483;
      ov(63 downto 0) := iv;
      ptr_deref_2507_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2507_root_address_inst
    process(ptr_deref_2507_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2507_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2507_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_2389_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2602_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2389_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2389_branch_req_0,
          ack0 => do_while_stmt_2389_branch_ack_0,
          ack1 => do_while_stmt_2389_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2603_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_2599;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2603_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2603_branch_req_0,
          ack0 => if_stmt_2603_branch_ack_0,
          ack1 => if_stmt_2603_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2309_inst
    process(call7_2251) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2251, type_cast_2308_wire_constant, tmp_var);
      add45_2310 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2320_inst
    process(call9_2254) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2254, type_cast_2319_wire_constant, tmp_var);
      add58_2321 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2339_inst
    process(call3_2245) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call3_2245, type_cast_2338_wire_constant, tmp_var);
      sub91_2340 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2425_inst
    process(sub_2315, mul_2421) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2315, mul_2421, tmp_var);
      sub48_2426 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2435_inst
    process(sub61_2326, mul54_2431) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2326, mul54_2431, tmp_var);
      sub62_2436 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2528_inst
    process(input_dim2x_x1_2396) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2396, type_cast_2527_wire_constant, tmp_var);
      add101_2529 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2556_inst
    process(inc_2549, input_dim1x_x1_2513_delayed_2_0_2552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc_2549, input_dim1x_x1_2513_delayed_2_0_2552, tmp_var);
      input_dim1x_x0_2557 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2573_inst
    process(inc113_2566, input_dim0x_x1_2527_delayed_3_0_2569) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc113_2566, input_dim0x_x1_2527_delayed_3_0_2569, tmp_var);
      inc113x_xinput_dim0x_x1_2574 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2365_inst
    process(shr120140_2355, shr124141_2361) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr120140_2355, shr124141_2361, tmp_var);
      add125_2366 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2415_inst
    process(add_2288, indvar_2391) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2288, indvar_2391, tmp_var);
      add_src_0x_x0_2416 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2595_inst
    process(indvar_2391) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2391, type_cast_2594_wire_constant, tmp_var);
      indvarx_xnext_2596 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2457_inst
    process(mul76_2453, conv70_2444) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2453, conv70_2444, tmp_var);
      add77_2458 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2467_inst
    process(mul78_2463, conv65_2440) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2463, conv65_2440, tmp_var);
      add79_2468 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2494_inst
    process(shr84_2489) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr84_2489, type_cast_2493_wire_constant, tmp_var);
      idxprom85_2495 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2561_inst
    process(input_dim1x_x0_2557, call1_2242) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1x_x0_2557, call1_2242, tmp_var);
      cmp109_2562 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2589_inst
    process(conv116_2585, add125_2366) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv116_2585, add125_2366, tmp_var);
      cmp126_2590 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2303_inst
    process(call_2239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2239, type_cast_2302_wire_constant, tmp_var);
      shr139_2304 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2354_inst
    process(conv119_2349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv119_2349, type_cast_2353_wire_constant, tmp_var);
      shr120140_2355 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2360_inst
    process(conv119_2349) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv119_2349, type_cast_2359_wire_constant, tmp_var);
      shr124141_2361 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2488_inst
    process(add79_2468) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2468, type_cast_2487_wire_constant, tmp_var);
      shr84_2489 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2420_inst
    process(input_dim0x_x1_2406, call13_2260) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x1_2406, call13_2260, tmp_var);
      mul_2421 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2430_inst
    process(input_dim1x_x1_2401, call13_2260) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2401, call13_2260, tmp_var);
      mul54_2431 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2452_inst
    process(conv75_2448, conv73_2334) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2448, conv73_2334, tmp_var);
      mul76_2453 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2462_inst
    process(add77_2458, conv68_2330) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2458, conv68_2330, tmp_var);
      mul78_2463 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2602_inst
    process(cmp126_2590) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp126_2590, tmp_var);
      NOT_u1_u1_2602_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u32_u32_2287_inst
    process(shl_2276, conv17_2283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2276, conv17_2283, tmp_var);
      add_2288 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2275_inst
    process(conv_2270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2270, type_cast_2274_wire_constant, tmp_var);
      shl_2276 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2522_inst
    process(type_cast_2520_wire, type_cast_2485_2485_delayed_2_0_2517) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2520_wire, type_cast_2485_2485_delayed_2_0_2517, tmp_var);
      cmp_2523 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2314_inst
    process(add45_2310, call14_2263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2310, call14_2263, tmp_var);
      sub_2315 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2325_inst
    process(add58_2321, call14_2263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2321, call14_2263, tmp_var);
      sub61_2326 <= tmp_var; --
    end process;
    -- binary operator XOR_u16_u16_2548_inst
    process(iNsTr_18_2543) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntXor_proc(iNsTr_18_2543, type_cast_2547_wire_constant, tmp_var);
      inc_2549 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2477_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2476_scaled;
      array_obj_ref_2477_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2477_index_offset_req_0;
      array_obj_ref_2477_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2477_index_offset_req_1;
      array_obj_ref_2477_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2500_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom85_2499_scaled;
      array_obj_ref_2500_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2500_index_offset_req_0;
      array_obj_ref_2500_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2500_index_offset_req_1;
      array_obj_ref_2500_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- unary operator type_cast_2343_inst
    process(sub91_2340) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", sub91_2340, tmp_var);
      type_cast_2343_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2482_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2482_load_0_req_0;
      ptr_deref_2482_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2482_load_0_req_1;
      ptr_deref_2482_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2482_word_address_0;
      ptr_deref_2482_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2507_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2507_store_0_req_0;
      ptr_deref_2507_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2507_store_0_req_1;
      ptr_deref_2507_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2507_word_address_0;
      data_in <= ptr_deref_2507_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2259_inst RPIPE_Block2_start_2278_inst RPIPE_Block2_start_2262_inst RPIPE_Block2_start_2265_inst RPIPE_Block2_start_2290_inst RPIPE_Block2_start_2293_inst RPIPE_Block2_start_2296_inst RPIPE_Block2_start_2256_inst RPIPE_Block2_start_2253_inst RPIPE_Block2_start_2250_inst RPIPE_Block2_start_2247_inst RPIPE_Block2_start_2244_inst RPIPE_Block2_start_2241_inst RPIPE_Block2_start_2238_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2259_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2278_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2262_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2265_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2290_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2293_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2296_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2256_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2253_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2250_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2247_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2244_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2241_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2238_inst_req_0;
      RPIPE_Block2_start_2259_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2278_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2262_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2265_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2290_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2293_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2296_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2256_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2253_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2250_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2247_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2244_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2241_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2238_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2259_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2278_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2262_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2265_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2290_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2293_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2296_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2256_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2253_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2250_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2247_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2244_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2241_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2238_inst_req_1;
      RPIPE_Block2_start_2259_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2278_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2262_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2265_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2290_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2293_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2296_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2256_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2253_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2250_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2247_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2244_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2241_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2238_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call13_2260 <= data_out(223 downto 208);
      call16_2279 <= data_out(207 downto 192);
      call14_2263 <= data_out(191 downto 176);
      call15_2266 <= data_out(175 downto 160);
      call18_2291 <= data_out(159 downto 144);
      call20_2294 <= data_out(143 downto 128);
      call22_2297 <= data_out(127 downto 112);
      call11_2257 <= data_out(111 downto 96);
      call9_2254 <= data_out(95 downto 80);
      call7_2251 <= data_out(79 downto 64);
      call5_2248 <= data_out(63 downto 48);
      call3_2245 <= data_out(47 downto 32);
      call1_2242 <= data_out(31 downto 16);
      call_2239 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2609_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2609_inst_req_0;
      WPIPE_Block2_done_2609_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2609_inst_req_1;
      WPIPE_Block2_done_2609_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2611_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6687_start: Boolean;
  signal convTransposeD_CP_6687_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2641_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2678_inst_ack_1 : boolean;
  signal type_cast_2726_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2623_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2626_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2678_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2635_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2660_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2660_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2675_inst_ack_0 : boolean;
  signal type_cast_2737_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2635_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2635_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2647_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2632_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2660_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2660_inst_ack_1 : boolean;
  signal type_cast_2737_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2626_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2647_inst_ack_0 : boolean;
  signal type_cast_2737_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2647_inst_req_1 : boolean;
  signal type_cast_2651_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2678_inst_req_0 : boolean;
  signal type_cast_2726_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2632_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2647_inst_ack_1 : boolean;
  signal type_cast_2651_inst_req_1 : boolean;
  signal do_while_stmt_2761_branch_req_0 : boolean;
  signal W_add106_2853_delayed_1_0_2902_inst_req_0 : boolean;
  signal type_cast_2664_inst_req_0 : boolean;
  signal type_cast_2664_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2675_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2641_inst_ack_0 : boolean;
  signal type_cast_2726_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2675_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2620_inst_req_0 : boolean;
  signal type_cast_2737_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2623_inst_req_1 : boolean;
  signal type_cast_2664_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2675_inst_ack_1 : boolean;
  signal type_cast_2664_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2635_inst_ack_0 : boolean;
  signal type_cast_2888_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2641_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2638_inst_ack_1 : boolean;
  signal type_cast_2888_inst_ack_1 : boolean;
  signal type_cast_2651_inst_req_0 : boolean;
  signal type_cast_2722_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2626_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2632_inst_req_1 : boolean;
  signal type_cast_2651_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2620_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2626_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2678_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2644_inst_req_0 : boolean;
  signal type_cast_2722_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2629_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2620_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2638_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2620_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2644_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2638_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2672_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2672_inst_ack_0 : boolean;
  signal type_cast_2726_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2638_inst_req_1 : boolean;
  signal type_cast_2722_inst_req_1 : boolean;
  signal W_add106_2853_delayed_1_0_2902_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2644_inst_ack_1 : boolean;
  signal W_input_dim0x_x1_2884_delayed_3_0_2939_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2644_inst_req_1 : boolean;
  signal do_while_stmt_2761_branch_ack_0 : boolean;
  signal type_cast_2888_inst_ack_0 : boolean;
  signal phi_stmt_2763_ack_0 : boolean;
  signal RPIPE_Block3_start_2632_inst_ack_1 : boolean;
  signal do_while_stmt_2761_branch_ack_1 : boolean;
  signal RPIPE_Block3_start_2672_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2672_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2623_inst_ack_0 : boolean;
  signal phi_stmt_2763_req_1 : boolean;
  signal RPIPE_Block3_start_2623_inst_req_0 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal type_cast_2766_inst_req_1 : boolean;
  signal type_cast_2766_inst_ack_1 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal type_cast_2888_inst_req_0 : boolean;
  signal phi_stmt_2763_req_0 : boolean;
  signal phi_stmt_2756_req_0 : boolean;
  signal type_cast_2759_inst_ack_1 : boolean;
  signal phi_stmt_2768_req_0 : boolean;
  signal phi_stmt_2768_req_1 : boolean;
  signal phi_stmt_2768_ack_0 : boolean;
  signal type_cast_2722_inst_ack_1 : boolean;
  signal type_cast_2884_inst_req_0 : boolean;
  signal type_cast_2759_inst_req_1 : boolean;
  signal type_cast_2771_inst_req_0 : boolean;
  signal type_cast_2771_inst_ack_0 : boolean;
  signal type_cast_2771_inst_req_1 : boolean;
  signal type_cast_2771_inst_ack_1 : boolean;
  signal W_input_dim0x_x1_2884_delayed_3_0_2939_inst_req_1 : boolean;
  signal W_input_dim0x_x1_2884_delayed_3_0_2939_inst_ack_0 : boolean;
  signal W_input_dim0x_x1_2884_delayed_3_0_2939_inst_req_0 : boolean;
  signal phi_stmt_2773_req_0 : boolean;
  signal phi_stmt_2773_req_1 : boolean;
  signal phi_stmt_2773_ack_0 : boolean;
  signal type_cast_2937_inst_ack_1 : boolean;
  signal type_cast_2776_inst_req_0 : boolean;
  signal type_cast_2759_inst_ack_0 : boolean;
  signal type_cast_2776_inst_ack_0 : boolean;
  signal type_cast_2776_inst_req_1 : boolean;
  signal type_cast_2759_inst_req_0 : boolean;
  signal type_cast_2776_inst_ack_1 : boolean;
  signal type_cast_2937_inst_req_1 : boolean;
  signal type_cast_2937_inst_ack_0 : boolean;
  signal phi_stmt_2778_req_0 : boolean;
  signal phi_stmt_2778_req_1 : boolean;
  signal phi_stmt_2778_ack_0 : boolean;
  signal type_cast_2937_inst_req_0 : boolean;
  signal type_cast_2781_inst_req_0 : boolean;
  signal type_cast_2781_inst_ack_0 : boolean;
  signal type_cast_2781_inst_req_1 : boolean;
  signal type_cast_2781_inst_ack_1 : boolean;
  signal input_dim0x_x1_at_entry_2756_2782_buf_req_0 : boolean;
  signal input_dim0x_x1_at_entry_2756_2782_buf_ack_0 : boolean;
  signal input_dim0x_x1_at_entry_2756_2782_buf_req_1 : boolean;
  signal input_dim0x_x1_at_entry_2756_2782_buf_ack_1 : boolean;
  signal type_cast_2811_inst_req_0 : boolean;
  signal type_cast_2811_inst_ack_0 : boolean;
  signal if_stmt_2971_branch_ack_0 : boolean;
  signal type_cast_2811_inst_req_1 : boolean;
  signal type_cast_2811_inst_ack_1 : boolean;
  signal type_cast_2815_inst_req_0 : boolean;
  signal type_cast_2815_inst_ack_0 : boolean;
  signal type_cast_2815_inst_req_1 : boolean;
  signal type_cast_2815_inst_ack_1 : boolean;
  signal W_input_dim1x_x1_2870_delayed_2_0_2922_inst_ack_1 : boolean;
  signal W_input_dim1x_x1_2870_delayed_2_0_2922_inst_req_1 : boolean;
  signal type_cast_2819_inst_req_0 : boolean;
  signal type_cast_2819_inst_ack_0 : boolean;
  signal type_cast_2819_inst_req_1 : boolean;
  signal type_cast_2819_inst_ack_1 : boolean;
  signal ptr_deref_2879_store_0_ack_1 : boolean;
  signal type_cast_2843_inst_req_0 : boolean;
  signal type_cast_2843_inst_ack_0 : boolean;
  signal if_stmt_2971_branch_ack_1 : boolean;
  signal type_cast_2843_inst_req_1 : boolean;
  signal type_cast_2843_inst_ack_1 : boolean;
  signal ptr_deref_2879_store_0_req_1 : boolean;
  signal W_input_dim1x_x1_2870_delayed_2_0_2922_inst_ack_0 : boolean;
  signal W_input_dim1x_x1_2870_delayed_2_0_2922_inst_req_0 : boolean;
  signal array_obj_ref_2849_index_offset_req_0 : boolean;
  signal WPIPE_Block3_done_2977_inst_ack_1 : boolean;
  signal array_obj_ref_2849_index_offset_ack_0 : boolean;
  signal array_obj_ref_2849_index_offset_req_1 : boolean;
  signal WPIPE_Block3_done_2977_inst_req_1 : boolean;
  signal array_obj_ref_2849_index_offset_ack_1 : boolean;
  signal addr_of_2850_final_reg_req_0 : boolean;
  signal WPIPE_Block3_done_2977_inst_ack_0 : boolean;
  signal addr_of_2850_final_reg_ack_0 : boolean;
  signal if_stmt_2971_branch_req_0 : boolean;
  signal addr_of_2850_final_reg_req_1 : boolean;
  signal WPIPE_Block3_done_2977_inst_req_0 : boolean;
  signal addr_of_2850_final_reg_ack_1 : boolean;
  signal ptr_deref_2854_load_0_req_0 : boolean;
  signal ptr_deref_2854_load_0_ack_0 : boolean;
  signal type_cast_2884_inst_ack_0 : boolean;
  signal ptr_deref_2854_load_0_req_1 : boolean;
  signal type_cast_2914_inst_ack_1 : boolean;
  signal ptr_deref_2854_load_0_ack_1 : boolean;
  signal type_cast_2914_inst_req_1 : boolean;
  signal type_cast_2884_inst_ack_1 : boolean;
  signal type_cast_2884_inst_req_1 : boolean;
  signal phi_stmt_2756_ack_0 : boolean;
  signal type_cast_2914_inst_ack_0 : boolean;
  signal type_cast_2914_inst_req_0 : boolean;
  signal W_add106_2853_delayed_1_0_2902_inst_ack_1 : boolean;
  signal W_add106_2853_delayed_1_0_2902_inst_req_1 : boolean;
  signal array_obj_ref_2872_index_offset_req_0 : boolean;
  signal array_obj_ref_2872_index_offset_ack_0 : boolean;
  signal array_obj_ref_2872_index_offset_req_1 : boolean;
  signal array_obj_ref_2872_index_offset_ack_1 : boolean;
  signal addr_of_2873_final_reg_req_0 : boolean;
  signal addr_of_2873_final_reg_ack_0 : boolean;
  signal addr_of_2873_final_reg_req_1 : boolean;
  signal addr_of_2873_final_reg_ack_1 : boolean;
  signal W_arrayidx91_2830_delayed_6_0_2875_inst_req_0 : boolean;
  signal W_arrayidx91_2830_delayed_6_0_2875_inst_ack_0 : boolean;
  signal W_arrayidx91_2830_delayed_6_0_2875_inst_req_1 : boolean;
  signal W_arrayidx91_2830_delayed_6_0_2875_inst_ack_1 : boolean;
  signal ptr_deref_2879_store_0_req_0 : boolean;
  signal ptr_deref_2879_store_0_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6687_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6687_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6687_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6687_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6687: Block -- control-path 
    signal convTransposeD_CP_6687_elements: BooleanArray(220 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6687_elements(0) <= convTransposeD_CP_6687_start;
    convTransposeD_CP_6687_symbol <= convTransposeD_CP_6687_elements(216);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2618/$entry
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/$entry
      -- CP-element group 0: 	 branch_block_stmt_2618/branch_block_stmt_2618__entry__
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679__entry__
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Update/cr
      -- 
    cr_6866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(0), ack => type_cast_2651_inst_req_1); -- 
    rr_6721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(0), ack => RPIPE_Block3_start_2620_inst_req_0); -- 
    cr_6894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(0), ack => type_cast_2664_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	212 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	213 
    -- CP-element group 1: 	214 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971__entry__
      -- CP-element group 1: 	 branch_block_stmt_2618/do_while_stmt_2761__exit__
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_2618/R_whilex_xbody_whilex_xend_taken_2972_place
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_2618/if_stmt_2971_eval_test/$exit
      -- 
    branch_req_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(1), ack => if_stmt_2971_branch_req_0); -- 
    convTransposeD_CP_6687_elements(1) <= convTransposeD_CP_6687_elements(212);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Update/cr
      -- 
    ra_6722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2620_inst_ack_0, ack => convTransposeD_CP_6687_elements(2)); -- 
    cr_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(2), ack => RPIPE_Block3_start_2620_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2620_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Sample/$entry
      -- 
    ca_6727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2620_inst_ack_1, ack => convTransposeD_CP_6687_elements(3)); -- 
    rr_6735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(3), ack => RPIPE_Block3_start_2623_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_sample_completed_
      -- 
    ra_6736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2623_inst_ack_0, ack => convTransposeD_CP_6687_elements(4)); -- 
    cr_6740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(4), ack => RPIPE_Block3_start_2623_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2623_update_completed_
      -- 
    ca_6741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2623_inst_ack_1, ack => convTransposeD_CP_6687_elements(5)); -- 
    rr_6749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(5), ack => RPIPE_Block3_start_2626_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Update/$entry
      -- 
    ra_6750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2626_inst_ack_0, ack => convTransposeD_CP_6687_elements(6)); -- 
    cr_6754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(6), ack => RPIPE_Block3_start_2626_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2626_update_completed_
      -- 
    ca_6755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2626_inst_ack_1, ack => convTransposeD_CP_6687_elements(7)); -- 
    rr_6763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(7), ack => RPIPE_Block3_start_2629_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Update/cr
      -- 
    ra_6764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2629_inst_ack_0, ack => convTransposeD_CP_6687_elements(8)); -- 
    cr_6768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(8), ack => RPIPE_Block3_start_2629_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2629_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_sample_start_
      -- 
    ca_6769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2629_inst_ack_1, ack => convTransposeD_CP_6687_elements(9)); -- 
    rr_6777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(9), ack => RPIPE_Block3_start_2632_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_sample_completed_
      -- 
    ra_6778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2632_inst_ack_0, ack => convTransposeD_CP_6687_elements(10)); -- 
    cr_6782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(10), ack => RPIPE_Block3_start_2632_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2632_Update/ca
      -- 
    ca_6783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2632_inst_ack_1, ack => convTransposeD_CP_6687_elements(11)); -- 
    rr_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(11), ack => RPIPE_Block3_start_2635_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_update_start_
      -- 
    ra_6792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2635_inst_ack_0, ack => convTransposeD_CP_6687_elements(12)); -- 
    cr_6796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(12), ack => RPIPE_Block3_start_2635_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2635_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Sample/rr
      -- 
    ca_6797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2635_inst_ack_1, ack => convTransposeD_CP_6687_elements(13)); -- 
    rr_6805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(13), ack => RPIPE_Block3_start_2638_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Update/cr
      -- 
    ra_6806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2638_inst_ack_0, ack => convTransposeD_CP_6687_elements(14)); -- 
    cr_6810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(14), ack => RPIPE_Block3_start_2638_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2638_Update/$exit
      -- 
    ca_6811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2638_inst_ack_1, ack => convTransposeD_CP_6687_elements(15)); -- 
    rr_6819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(15), ack => RPIPE_Block3_start_2641_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_sample_completed_
      -- 
    ra_6820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2641_inst_ack_0, ack => convTransposeD_CP_6687_elements(16)); -- 
    cr_6824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(16), ack => RPIPE_Block3_start_2641_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2641_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Sample/rr
      -- 
    ca_6825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2641_inst_ack_1, ack => convTransposeD_CP_6687_elements(17)); -- 
    rr_6833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(17), ack => RPIPE_Block3_start_2644_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Update/$entry
      -- 
    ra_6834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2644_inst_ack_0, ack => convTransposeD_CP_6687_elements(18)); -- 
    cr_6838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(18), ack => RPIPE_Block3_start_2644_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2644_Update/$exit
      -- 
    ca_6839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2644_inst_ack_1, ack => convTransposeD_CP_6687_elements(19)); -- 
    rr_6847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(19), ack => RPIPE_Block3_start_2647_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Sample/$exit
      -- 
    ra_6848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2647_inst_ack_0, ack => convTransposeD_CP_6687_elements(20)); -- 
    cr_6852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(20), ack => RPIPE_Block3_start_2647_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2647_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Sample/rr
      -- 
    ca_6853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2647_inst_ack_1, ack => convTransposeD_CP_6687_elements(21)); -- 
    rr_6861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(21), ack => type_cast_2651_inst_req_0); -- 
    rr_6875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(21), ack => RPIPE_Block3_start_2660_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Sample/ra
      -- 
    ra_6862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2651_inst_ack_0, ack => convTransposeD_CP_6687_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2651_Update/$exit
      -- 
    ca_6867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2651_inst_ack_1, ack => convTransposeD_CP_6687_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_update_start_
      -- 
    ra_6876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2660_inst_ack_0, ack => convTransposeD_CP_6687_elements(24)); -- 
    cr_6880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(24), ack => RPIPE_Block3_start_2660_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2660_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Sample/rr
      -- 
    ca_6881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2660_inst_ack_1, ack => convTransposeD_CP_6687_elements(25)); -- 
    rr_6889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(25), ack => type_cast_2664_inst_req_0); -- 
    rr_6903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(25), ack => RPIPE_Block3_start_2672_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Sample/ra
      -- 
    ra_6890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2664_inst_ack_0, ack => convTransposeD_CP_6687_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/type_cast_2664_Update/ca
      -- 
    ca_6895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2664_inst_ack_1, ack => convTransposeD_CP_6687_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Update/cr
      -- 
    ra_6904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2672_inst_ack_0, ack => convTransposeD_CP_6687_elements(28)); -- 
    cr_6908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(28), ack => RPIPE_Block3_start_2672_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2672_Update/$exit
      -- 
    ca_6909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2672_inst_ack_1, ack => convTransposeD_CP_6687_elements(29)); -- 
    rr_6917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(29), ack => RPIPE_Block3_start_2675_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_sample_completed_
      -- 
    ra_6918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2675_inst_ack_0, ack => convTransposeD_CP_6687_elements(30)); -- 
    cr_6922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(30), ack => RPIPE_Block3_start_2675_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2675_update_completed_
      -- 
    ca_6923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2675_inst_ack_1, ack => convTransposeD_CP_6687_elements(31)); -- 
    rr_6931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(31), ack => RPIPE_Block3_start_2678_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Update/$entry
      -- 
    ra_6932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2678_inst_ack_0, ack => convTransposeD_CP_6687_elements(32)); -- 
    cr_6936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(32), ack => RPIPE_Block3_start_2678_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/RPIPE_Block3_start_2678_Update/$exit
      -- 
    ca_6937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2678_inst_ack_1, ack => convTransposeD_CP_6687_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679/$exit
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2621_to_assign_stmt_2679__exit__
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738__entry__
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_sample_start_
      -- 
    cr_6981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(34), ack => type_cast_2737_inst_req_1); -- 
    rr_6962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(34), ack => type_cast_2726_inst_req_0); -- 
    rr_6976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(34), ack => type_cast_2737_inst_req_0); -- 
    rr_6948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(34), ack => type_cast_2722_inst_req_0); -- 
    cr_6967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(34), ack => type_cast_2726_inst_req_1); -- 
    cr_6953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(34), ack => type_cast_2722_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(23) & convTransposeD_CP_6687_elements(27) & convTransposeD_CP_6687_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Sample/ra
      -- 
    ra_6949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_0, ack => convTransposeD_CP_6687_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2722_Update/ca
      -- 
    ca_6954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_1, ack => convTransposeD_CP_6687_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_sample_completed_
      -- 
    ra_6963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_0, ack => convTransposeD_CP_6687_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2726_update_completed_
      -- 
    ca_6968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_1, ack => convTransposeD_CP_6687_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_sample_completed_
      -- 
    ra_6977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2737_inst_ack_0, ack => convTransposeD_CP_6687_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/type_cast_2737_update_completed_
      -- 
    ca_6982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2737_inst_ack_1, ack => convTransposeD_CP_6687_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	217 
    -- CP-element group 41: 	218 
    -- CP-element group 41:  members (12) 
      -- CP-element group 41: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738/$exit
      -- CP-element group 41: 	 branch_block_stmt_2618/assign_stmt_2686_to_assign_stmt_2738__exit__
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/cr
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/$entry
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/$entry
      -- CP-element group 41: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/$entry
      -- 
    cr_7617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(41), ack => type_cast_2759_inst_req_1); -- 
    rr_7612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(41), ack => type_cast_2759_inst_req_0); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(36) & convTransposeD_CP_6687_elements(38) & convTransposeD_CP_6687_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  place  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	220 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	48 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761__entry__
      -- CP-element group 42: 	 branch_block_stmt_2618/do_while_stmt_2761/$entry
      -- 
    convTransposeD_CP_6687_elements(42) <= convTransposeD_CP_6687_elements(220);
    -- CP-element group 43:  merge  place  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	212 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761__exit__
      -- 
    -- Element group convTransposeD_CP_6687_elements(43) is bound as output of CP function.
    -- CP-element group 44:  merge  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_back
      -- 
    -- Element group convTransposeD_CP_6687_elements(44) is bound as output of CP function.
    -- CP-element group 45:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	50 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	210 
    -- CP-element group 45: 	211 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2618/do_while_stmt_2761/condition_done
      -- CP-element group 45: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_taken/$entry
      -- CP-element group 45: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_exit/$entry
      -- 
    convTransposeD_CP_6687_elements(45) <= convTransposeD_CP_6687_elements(50);
    -- CP-element group 46:  branch  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	209 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_body_done
      -- 
    convTransposeD_CP_6687_elements(46) <= convTransposeD_CP_6687_elements(209);
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	59 
    -- CP-element group 47: 	80 
    -- CP-element group 47: 	101 
    -- CP-element group 47: 	122 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/back_edge_to_loop_body
      -- 
    convTransposeD_CP_6687_elements(47) <= convTransposeD_CP_6687_elements(44);
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	42 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	61 
    -- CP-element group 48: 	82 
    -- CP-element group 48: 	103 
    -- CP-element group 48: 	124 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/first_time_through_loop_body
      -- 
    convTransposeD_CP_6687_elements(48) <= convTransposeD_CP_6687_elements(42);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	55 
    -- CP-element group 49: 	56 
    -- CP-element group 49: 	74 
    -- CP-element group 49: 	75 
    -- CP-element group 49: 	95 
    -- CP-element group 49: 	96 
    -- CP-element group 49: 	116 
    -- CP-element group 49: 	117 
    -- CP-element group 49: 	154 
    -- CP-element group 49: 	155 
    -- CP-element group 49: 	165 
    -- CP-element group 49: 	167 
    -- CP-element group 49: 	184 
    -- CP-element group 49: 	208 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/$entry
      -- CP-element group 49: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/loop_body_start
      -- 
    -- Element group convTransposeD_CP_6687_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	54 
    -- CP-element group 50: 	203 
    -- CP-element group 50: 	207 
    -- CP-element group 50: 	208 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	45 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/condition_evaluated
      -- 
    condition_evaluated_6997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(50), ack => do_while_stmt_2761_branch_req_0); -- 
    convTransposeD_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(54) & convTransposeD_CP_6687_elements(203) & convTransposeD_CP_6687_elements(207) & convTransposeD_CP_6687_elements(208);
      gj_convTransposeD_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	55 
    -- CP-element group 51: 	74 
    -- CP-element group 51: 	95 
    -- CP-element group 51: 	116 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	76 
    -- CP-element group 51: 	97 
    -- CP-element group 51: 	118 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/aggregated_phi_sample_req
      -- 
    convTransposeD_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(55) & convTransposeD_CP_6687_elements(74) & convTransposeD_CP_6687_elements(95) & convTransposeD_CP_6687_elements(116) & convTransposeD_CP_6687_elements(54);
      gj_convTransposeD_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	57 
    -- CP-element group 52: 	77 
    -- CP-element group 52: 	98 
    -- CP-element group 52: 	119 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	181 
    -- CP-element group 52: 	185 
    -- CP-element group 52: 	189 
    -- CP-element group 52: 	193 
    -- CP-element group 52: 	197 
    -- CP-element group 52: 	201 
    -- CP-element group 52: 	205 
    -- CP-element group 52: 	209 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	55 
    -- CP-element group 52: 	74 
    -- CP-element group 52: 	95 
    -- CP-element group 52: 	116 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/aggregated_phi_sample_ack
      -- CP-element group 52: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_sample_completed_
      -- 
    convTransposeD_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(57) & convTransposeD_CP_6687_elements(77) & convTransposeD_CP_6687_elements(98) & convTransposeD_CP_6687_elements(119);
      gj_convTransposeD_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: 	75 
    -- CP-element group 53: 	96 
    -- CP-element group 53: 	117 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53: 	99 
    -- CP-element group 53: 	120 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/aggregated_phi_update_req
      -- 
    convTransposeD_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(56) & convTransposeD_CP_6687_elements(75) & convTransposeD_CP_6687_elements(96) & convTransposeD_CP_6687_elements(117);
      gj_convTransposeD_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	58 
    -- CP-element group 54: 	79 
    -- CP-element group 54: 	100 
    -- CP-element group 54: 	121 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	50 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/aggregated_phi_update_ack
      -- 
    convTransposeD_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(58) & convTransposeD_CP_6687_elements(79) & convTransposeD_CP_6687_elements(100) & convTransposeD_CP_6687_elements(121);
      gj_convTransposeD_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	49 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	51 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_sample_start_
      -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(52);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	49 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	151 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_update_start_
      -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(58) & convTransposeD_CP_6687_elements(151);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	52 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_sample_completed__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(57) is bound as output of CP function.
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	54 
    -- CP-element group 58: 	149 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_update_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	47 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_loopback_trigger
      -- 
    convTransposeD_CP_6687_elements(59) <= convTransposeD_CP_6687_elements(47);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_loopback_sample_req
      -- CP-element group 60: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_loopback_sample_req_ps
      -- 
    phi_stmt_2763_loopback_sample_req_7012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2763_loopback_sample_req_7012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(60), ack => phi_stmt_2763_req_0); -- 
    -- Element group convTransposeD_CP_6687_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	48 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_entry_trigger
      -- 
    convTransposeD_CP_6687_elements(61) <= convTransposeD_CP_6687_elements(48);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_entry_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_entry_sample_req
      -- 
    phi_stmt_2763_entry_sample_req_7015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2763_entry_sample_req_7015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(62), ack => phi_stmt_2763_req_1); -- 
    -- Element group convTransposeD_CP_6687_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_phi_mux_ack
      -- CP-element group 63: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2763_phi_mux_ack_ps
      -- 
    phi_stmt_2763_phi_mux_ack_7018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2763_ack_0, ack => convTransposeD_CP_6687_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_sample_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_update_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Sample/rr
      -- 
    rr_7031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(66), ack => type_cast_2766_inst_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(64) & convTransposeD_CP_6687_elements(68);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_update_start_
      -- CP-element group 67: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Update/$entry
      -- 
    cr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(67), ack => type_cast_2766_inst_req_1); -- 
    convTransposeD_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(65) & convTransposeD_CP_6687_elements(69);
      gj_convTransposeD_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Sample/ra
      -- 
    ra_7032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => convTransposeD_CP_6687_elements(68)); -- 
    -- CP-element group 69:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2766_Update/$exit
      -- 
    ca_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_1, ack => convTransposeD_CP_6687_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_sample_start__ps
      -- CP-element group 70: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_sample_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_update_start_
      -- CP-element group 71: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_update_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_update_completed__ps
      -- 
    convTransposeD_CP_6687_elements(72) <= convTransposeD_CP_6687_elements(73);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	72 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_indvar_at_entry_2767_update_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeD_CP_6687_elements(71), ack => convTransposeD_CP_6687_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	49 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	183 
    -- CP-element group 74: 	187 
    -- CP-element group 74: 	191 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	51 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_sample_start_
      -- 
    convTransposeD_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(183) & convTransposeD_CP_6687_elements(187) & convTransposeD_CP_6687_elements(191);
      gj_convTransposeD_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	49 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	139 
    -- CP-element group 75: 	182 
    -- CP-element group 75: 	190 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	53 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_update_start_
      -- 
    convTransposeD_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(79) & convTransposeD_CP_6687_elements(139) & convTransposeD_CP_6687_elements(182) & convTransposeD_CP_6687_elements(190);
      gj_convTransposeD_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	51 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_sample_start__ps
      -- 
    convTransposeD_CP_6687_elements(76) <= convTransposeD_CP_6687_elements(51);
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	52 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_sample_completed__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	53 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_update_start__ps
      -- 
    convTransposeD_CP_6687_elements(78) <= convTransposeD_CP_6687_elements(53);
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	54 
    -- CP-element group 79: 	137 
    -- CP-element group 79: 	180 
    -- CP-element group 79: 	188 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	75 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_update_completed__ps
      -- CP-element group 79: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_update_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	47 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_loopback_trigger
      -- 
    convTransposeD_CP_6687_elements(80) <= convTransposeD_CP_6687_elements(47);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_loopback_sample_req
      -- CP-element group 81: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_loopback_sample_req_ps
      -- 
    phi_stmt_2768_loopback_sample_req_7056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2768_loopback_sample_req_7056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(81), ack => phi_stmt_2768_req_0); -- 
    -- Element group convTransposeD_CP_6687_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	48 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_entry_trigger
      -- 
    convTransposeD_CP_6687_elements(82) <= convTransposeD_CP_6687_elements(48);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_entry_sample_req
      -- CP-element group 83: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_entry_sample_req_ps
      -- 
    phi_stmt_2768_entry_sample_req_7059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2768_entry_sample_req_7059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(83), ack => phi_stmt_2768_req_1); -- 
    -- Element group convTransposeD_CP_6687_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_phi_mux_ack
      -- CP-element group 84: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2768_phi_mux_ack_ps
      -- 
    phi_stmt_2768_phi_mux_ack_7062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2768_ack_0, ack => convTransposeD_CP_6687_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_sample_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_update_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Sample/rr
      -- 
    rr_7075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(87), ack => type_cast_2771_inst_req_0); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(85) & convTransposeD_CP_6687_elements(89);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_update_start_
      -- CP-element group 88: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Update/cr
      -- 
    cr_7080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(88), ack => type_cast_2771_inst_req_1); -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(86) & convTransposeD_CP_6687_elements(90);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Sample/ra
      -- 
    ra_7076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_0, ack => convTransposeD_CP_6687_elements(89)); -- 
    -- CP-element group 90:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2771_Update/ca
      -- 
    ca_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_1, ack => convTransposeD_CP_6687_elements(90)); -- 
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_sample_start__ps
      -- CP-element group 91: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_sample_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_update_start__ps
      -- CP-element group 92: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_update_start_
      -- 
    -- Element group convTransposeD_CP_6687_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_update_completed__ps
      -- 
    convTransposeD_CP_6687_elements(93) <= convTransposeD_CP_6687_elements(94);
    -- CP-element group 94:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	93 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim2x_x1_at_entry_2772_update_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(94) is a control-delay.
    cp_element_94_delay: control_delay_element  generic map(name => " 94_delay", delay_value => 1)  port map(req => convTransposeD_CP_6687_elements(92), ack => convTransposeD_CP_6687_elements(94), clk => clk, reset =>reset);
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	49 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	52 
    -- CP-element group 95: 	195 
    -- CP-element group 95: 	199 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	51 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_sample_start_
      -- 
    convTransposeD_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(195) & convTransposeD_CP_6687_elements(199);
      gj_convTransposeD_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	49 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	100 
    -- CP-element group 96: 	143 
    -- CP-element group 96: 	198 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	53 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_update_start_
      -- 
    convTransposeD_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(100) & convTransposeD_CP_6687_elements(143) & convTransposeD_CP_6687_elements(198);
      gj_convTransposeD_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	51 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_sample_start__ps
      -- 
    convTransposeD_CP_6687_elements(97) <= convTransposeD_CP_6687_elements(51);
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	52 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_sample_completed__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	53 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_update_start__ps
      -- 
    convTransposeD_CP_6687_elements(99) <= convTransposeD_CP_6687_elements(53);
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	54 
    -- CP-element group 100: 	141 
    -- CP-element group 100: 	196 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	96 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_update_completed__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	47 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_loopback_trigger
      -- 
    convTransposeD_CP_6687_elements(101) <= convTransposeD_CP_6687_elements(47);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_loopback_sample_req
      -- CP-element group 102: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_loopback_sample_req_ps
      -- 
    phi_stmt_2773_loopback_sample_req_7100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2773_loopback_sample_req_7100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(102), ack => phi_stmt_2773_req_0); -- 
    -- Element group convTransposeD_CP_6687_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	48 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_entry_trigger
      -- 
    convTransposeD_CP_6687_elements(103) <= convTransposeD_CP_6687_elements(48);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_entry_sample_req
      -- CP-element group 104: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_entry_sample_req_ps
      -- 
    phi_stmt_2773_entry_sample_req_7103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2773_entry_sample_req_7103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(104), ack => phi_stmt_2773_req_1); -- 
    -- Element group convTransposeD_CP_6687_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_phi_mux_ack
      -- CP-element group 105: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2773_phi_mux_ack_ps
      -- 
    phi_stmt_2773_phi_mux_ack_7106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2773_ack_0, ack => convTransposeD_CP_6687_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_sample_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_update_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Sample/rr
      -- 
    rr_7119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(108), ack => type_cast_2776_inst_req_0); -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(106) & convTransposeD_CP_6687_elements(110);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_update_start_
      -- CP-element group 109: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Update/cr
      -- 
    cr_7124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(109), ack => type_cast_2776_inst_req_1); -- 
    convTransposeD_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(107) & convTransposeD_CP_6687_elements(111);
      gj_convTransposeD_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_sample_completed__ps
      -- CP-element group 110: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Sample/ra
      -- 
    ra_7120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2776_inst_ack_0, ack => convTransposeD_CP_6687_elements(110)); -- 
    -- CP-element group 111:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_update_completed__ps
      -- CP-element group 111: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2776_Update/ca
      -- 
    ca_7125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2776_inst_ack_1, ack => convTransposeD_CP_6687_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_sample_start__ps
      -- CP-element group 112: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_sample_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_update_start__ps
      -- CP-element group 113: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_update_start_
      -- 
    -- Element group convTransposeD_CP_6687_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_update_completed__ps
      -- 
    convTransposeD_CP_6687_elements(114) <= convTransposeD_CP_6687_elements(115);
    -- CP-element group 115:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	114 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim1x_x1_at_entry_2777_update_completed_
      -- 
    -- Element group convTransposeD_CP_6687_elements(115) is a control-delay.
    cp_element_115_delay: control_delay_element  generic map(name => " 115_delay", delay_value => 1)  port map(req => convTransposeD_CP_6687_elements(113), ack => convTransposeD_CP_6687_elements(115), clk => clk, reset =>reset);
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	49 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	52 
    -- CP-element group 116: 	203 
    -- CP-element group 116: 	207 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	51 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_sample_start_
      -- 
    convTransposeD_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(203) & convTransposeD_CP_6687_elements(207);
      gj_convTransposeD_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	49 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: 	147 
    -- CP-element group 117: 	206 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	53 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_update_start_
      -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(121) & convTransposeD_CP_6687_elements(147) & convTransposeD_CP_6687_elements(206);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	51 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_sample_start__ps
      -- 
    convTransposeD_CP_6687_elements(118) <= convTransposeD_CP_6687_elements(51);
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	52 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_sample_completed__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	53 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_update_start__ps
      -- 
    convTransposeD_CP_6687_elements(120) <= convTransposeD_CP_6687_elements(53);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	54 
    -- CP-element group 121: 	145 
    -- CP-element group 121: 	204 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_update_completed__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	47 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_loopback_trigger
      -- 
    convTransposeD_CP_6687_elements(122) <= convTransposeD_CP_6687_elements(47);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_loopback_sample_req_ps
      -- 
    phi_stmt_2778_loopback_sample_req_7144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2778_loopback_sample_req_7144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(123), ack => phi_stmt_2778_req_0); -- 
    -- Element group convTransposeD_CP_6687_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	48 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_entry_trigger
      -- 
    convTransposeD_CP_6687_elements(124) <= convTransposeD_CP_6687_elements(48);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_entry_sample_req_ps
      -- 
    phi_stmt_2778_entry_sample_req_7147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2778_entry_sample_req_7147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(125), ack => phi_stmt_2778_req_1); -- 
    -- Element group convTransposeD_CP_6687_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_phi_mux_ack_ps
      -- CP-element group 126: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/phi_stmt_2778_phi_mux_ack
      -- 
    phi_stmt_2778_phi_mux_ack_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2778_ack_0, ack => convTransposeD_CP_6687_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_sample_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_update_start__ps
      -- 
    -- Element group convTransposeD_CP_6687_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Sample/rr
      -- 
    rr_7163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(129), ack => type_cast_2781_inst_req_0); -- 
    convTransposeD_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(127) & convTransposeD_CP_6687_elements(131);
      gj_convTransposeD_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_update_start_
      -- CP-element group 130: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Update/cr
      -- 
    cr_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(130), ack => type_cast_2781_inst_req_1); -- 
    convTransposeD_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(128) & convTransposeD_CP_6687_elements(132);
      gj_convTransposeD_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_sample_completed__ps
      -- CP-element group 131: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Sample/ra
      -- 
    ra_7164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2781_inst_ack_0, ack => convTransposeD_CP_6687_elements(131)); -- 
    -- CP-element group 132:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_update_completed__ps
      -- CP-element group 132: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2781_Update/ca
      -- 
    ca_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2781_inst_ack_1, ack => convTransposeD_CP_6687_elements(132)); -- 
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Sample/req
      -- 
    req_7181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(133), ack => input_dim0x_x1_at_entry_2756_2782_buf_req_0); -- 
    -- Element group convTransposeD_CP_6687_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_update_start_
      -- CP-element group 134: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Update/req
      -- 
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(134), ack => input_dim0x_x1_at_entry_2756_2782_buf_req_1); -- 
    -- Element group convTransposeD_CP_6687_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Sample/ack
      -- 
    ack_7182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_dim0x_x1_at_entry_2756_2782_buf_ack_0, ack => convTransposeD_CP_6687_elements(135)); -- 
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_update_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/R_input_dim0x_x1_at_entry_2782_Update/ack
      -- 
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_dim0x_x1_at_entry_2756_2782_buf_ack_1, ack => convTransposeD_CP_6687_elements(136)); -- 
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	79 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Sample/rr
      -- 
    rr_7196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(137), ack => type_cast_2811_inst_req_0); -- 
    convTransposeD_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(79) & convTransposeD_CP_6687_elements(139);
      gj_convTransposeD_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: 	168 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_update_start_
      -- CP-element group 138: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Update/cr
      -- 
    cr_7201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(138), ack => type_cast_2811_inst_req_1); -- 
    convTransposeD_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(140) & convTransposeD_CP_6687_elements(168);
      gj_convTransposeD_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	75 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Sample/ra
      -- 
    ra_7197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2811_inst_ack_0, ack => convTransposeD_CP_6687_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	166 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2811_Update/ca
      -- 
    ca_7202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2811_inst_ack_1, ack => convTransposeD_CP_6687_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	100 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Sample/rr
      -- 
    rr_7210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(141), ack => type_cast_2815_inst_req_0); -- 
    convTransposeD_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(100) & convTransposeD_CP_6687_elements(143);
      gj_convTransposeD_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: 	168 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_update_start_
      -- CP-element group 142: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Update/cr
      -- 
    cr_7215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(142), ack => type_cast_2815_inst_req_1); -- 
    convTransposeD_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(144) & convTransposeD_CP_6687_elements(168);
      gj_convTransposeD_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	96 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Sample/ra
      -- 
    ra_7211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2815_inst_ack_0, ack => convTransposeD_CP_6687_elements(143)); -- 
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	166 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	142 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2815_Update/ca
      -- 
    ca_7216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2815_inst_ack_1, ack => convTransposeD_CP_6687_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	121 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Sample/rr
      -- 
    rr_7224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(145), ack => type_cast_2819_inst_req_0); -- 
    convTransposeD_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(121) & convTransposeD_CP_6687_elements(147);
      gj_convTransposeD_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: 	168 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_update_start_
      -- CP-element group 146: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Update/cr
      -- 
    cr_7229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(146), ack => type_cast_2819_inst_req_1); -- 
    convTransposeD_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(148) & convTransposeD_CP_6687_elements(168);
      gj_convTransposeD_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	117 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Sample/ra
      -- 
    ra_7225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2819_inst_ack_0, ack => convTransposeD_CP_6687_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	166 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2819_Update/ca
      -- 
    ca_7230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2819_inst_ack_1, ack => convTransposeD_CP_6687_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	58 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Sample/rr
      -- 
    rr_7238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(149), ack => type_cast_2843_inst_req_0); -- 
    convTransposeD_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(58) & convTransposeD_CP_6687_elements(151);
      gj_convTransposeD_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: 	156 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_update_start_
      -- CP-element group 150: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Update/cr
      -- 
    cr_7243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(150), ack => type_cast_2843_inst_req_1); -- 
    convTransposeD_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(152) & convTransposeD_CP_6687_elements(156);
      gj_convTransposeD_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	56 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Sample/ra
      -- 
    ra_7239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2843_inst_ack_0, ack => convTransposeD_CP_6687_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	156 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (16) 
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2843_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_resized_1
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_scaled_1
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_computed_1
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_resize_1/$entry
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_resize_1/$exit
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_resize_1/index_resize_req
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_resize_1/index_resize_ack
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_scale_1/$entry
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_scale_1/$exit
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_scale_1/scale_rename_req
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_index_scale_1/scale_rename_ack
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Sample/req
      -- 
    ca_7244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2843_inst_ack_1, ack => convTransposeD_CP_6687_elements(152)); -- 
    req_7269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(152), ack => array_obj_ref_2849_index_offset_req_0); -- 
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	157 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	158 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	158 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_request/$entry
      -- CP-element group 153: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_request/req
      -- 
    req_7284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(153), ack => addr_of_2850_final_reg_req_0); -- 
    convTransposeD_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(157) & convTransposeD_CP_6687_elements(158);
      gj_convTransposeD_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	49 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	159 
    -- CP-element group 154: 	162 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	159 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_update_start_
      -- CP-element group 154: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_complete/$entry
      -- CP-element group 154: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_complete/req
      -- 
    req_7289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(154), ack => addr_of_2850_final_reg_req_1); -- 
    convTransposeD_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(159) & convTransposeD_CP_6687_elements(162);
      gj_convTransposeD_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	49 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	158 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_update_start
      -- CP-element group 155: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Update/req
      -- 
    req_7274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(155), ack => array_obj_ref_2849_index_offset_req_1); -- 
    convTransposeD_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(157) & convTransposeD_CP_6687_elements(158);
      gj_convTransposeD_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	152 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	209 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	150 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_sample_complete
      -- CP-element group 156: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Sample/ack
      -- 
    ack_7270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2849_index_offset_ack_0, ack => convTransposeD_CP_6687_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	153 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (8) 
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_root_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_offset_calculated
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_final_index_sum_regn_Update/ack
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_base_plus_offset/$entry
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_base_plus_offset/$exit
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_base_plus_offset/sum_rename_req
      -- CP-element group 157: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2849_base_plus_offset/sum_rename_ack
      -- 
    ack_7275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2849_index_offset_ack_1, ack => convTransposeD_CP_6687_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	153 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	155 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_request/$exit
      -- CP-element group 158: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_request/ack
      -- 
    ack_7285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2850_final_reg_ack_0, ack => convTransposeD_CP_6687_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	154 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	154 
    -- CP-element group 159:  members (19) 
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_complete/$exit
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2850_complete/ack
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_word_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_root_address_calculated
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_address_resized
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_addr_resize/$entry
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_addr_resize/$exit
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_addr_resize/base_resize_req
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_addr_resize/base_resize_ack
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_plus_offset/$entry
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_plus_offset/$exit
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_plus_offset/sum_rename_req
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_base_plus_offset/sum_rename_ack
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_word_addrgen/$entry
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_word_addrgen/$exit
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_word_addrgen/root_register_req
      -- CP-element group 159: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_word_addrgen/root_register_ack
      -- 
    ack_7290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2850_final_reg_ack_1, ack => convTransposeD_CP_6687_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (5) 
      -- CP-element group 160: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/word_access_start/$entry
      -- CP-element group 160: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/word_access_start/word_0/$entry
      -- CP-element group 160: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/word_access_start/word_0/rr
      -- 
    rr_7323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(160), ack => ptr_deref_2854_load_0_req_0); -- 
    convTransposeD_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(159) & convTransposeD_CP_6687_elements(162);
      gj_convTransposeD_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	178 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_update_start_
      -- CP-element group 161: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/word_access_complete/$entry
      -- CP-element group 161: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/word_access_complete/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/word_access_complete/word_0/cr
      -- 
    cr_7334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(161), ack => ptr_deref_2854_load_0_req_1); -- 
    convTransposeD_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(163) & convTransposeD_CP_6687_elements(178);
      gj_convTransposeD_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	154 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Sample/word_access_start/word_0/ra
      -- 
    ra_7324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2854_load_0_ack_0, ack => convTransposeD_CP_6687_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	176 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/ptr_deref_2854_Merge/$entry
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/ptr_deref_2854_Merge/$exit
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/ptr_deref_2854_Merge/merge_req
      -- CP-element group 163: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2854_Update/ptr_deref_2854_Merge/merge_ack
      -- 
    ca_7335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2854_load_0_ack_1, ack => convTransposeD_CP_6687_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	169 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	170 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	170 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_request/$entry
      -- CP-element group 164: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_request/req
      -- 
    req_7380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(164), ack => addr_of_2873_final_reg_req_0); -- 
    convTransposeD_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(169) & convTransposeD_CP_6687_elements(170);
      gj_convTransposeD_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	49 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	171 
    -- CP-element group 165: 	174 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	171 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_update_start_
      -- CP-element group 165: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_complete/$entry
      -- CP-element group 165: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_complete/req
      -- 
    req_7385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(165), ack => addr_of_2873_final_reg_req_1); -- 
    convTransposeD_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(171) & convTransposeD_CP_6687_elements(174);
      gj_convTransposeD_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	140 
    -- CP-element group 166: 	144 
    -- CP-element group 166: 	148 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (13) 
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_resized_1
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_scaled_1
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_computed_1
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_resize_1/$entry
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_resize_1/$exit
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_resize_1/index_resize_req
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_resize_1/index_resize_ack
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_scale_1/$entry
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_scale_1/$exit
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_scale_1/scale_rename_req
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_index_scale_1/scale_rename_ack
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Sample/req
      -- 
    req_7365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(166), ack => array_obj_ref_2872_index_offset_req_0); -- 
    convTransposeD_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(140) & convTransposeD_CP_6687_elements(144) & convTransposeD_CP_6687_elements(148);
      gj_convTransposeD_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	49 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: 	170 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_update_start
      -- CP-element group 167: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Update/req
      -- 
    req_7370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(167), ack => array_obj_ref_2872_index_offset_req_1); -- 
    convTransposeD_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(169) & convTransposeD_CP_6687_elements(170);
      gj_convTransposeD_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	209 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	138 
    -- CP-element group 168: 	142 
    -- CP-element group 168: 	146 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_sample_complete
      -- CP-element group 168: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Sample/ack
      -- 
    ack_7366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2872_index_offset_ack_0, ack => convTransposeD_CP_6687_elements(168)); -- 
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	164 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (8) 
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_root_address_calculated
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_offset_calculated
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_final_index_sum_regn_Update/ack
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_base_plus_offset/$entry
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_base_plus_offset/$exit
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_base_plus_offset/sum_rename_req
      -- CP-element group 169: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/array_obj_ref_2872_base_plus_offset/sum_rename_ack
      -- 
    ack_7371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2872_index_offset_ack_1, ack => convTransposeD_CP_6687_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	164 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	164 
    -- CP-element group 170: 	167 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_request/$exit
      -- CP-element group 170: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_request/ack
      -- 
    ack_7381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2873_final_reg_ack_0, ack => convTransposeD_CP_6687_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	165 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	165 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_complete/$exit
      -- CP-element group 171: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/addr_of_2873_complete/ack
      -- 
    ack_7386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2873_final_reg_ack_1, ack => convTransposeD_CP_6687_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Sample/req
      -- 
    req_7394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(172), ack => W_arrayidx91_2830_delayed_6_0_2875_inst_req_0); -- 
    convTransposeD_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(171) & convTransposeD_CP_6687_elements(174);
      gj_convTransposeD_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	178 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_update_start_
      -- CP-element group 173: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Update/req
      -- 
    req_7399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(173), ack => W_arrayidx91_2830_delayed_6_0_2875_inst_req_1); -- 
    convTransposeD_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(175) & convTransposeD_CP_6687_elements(178);
      gj_convTransposeD_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	165 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Sample/ack
      -- 
    ack_7395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx91_2830_delayed_6_0_2875_inst_ack_0, ack => convTransposeD_CP_6687_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (19) 
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2877_Update/ack
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_address_calculated
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_word_address_calculated
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_root_address_calculated
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_address_resized
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_addr_resize/$entry
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_addr_resize/$exit
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_addr_resize/base_resize_req
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_addr_resize/base_resize_ack
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_plus_offset/$entry
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_plus_offset/$exit
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_plus_offset/sum_rename_req
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_base_plus_offset/sum_rename_ack
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_word_addrgen/$entry
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_word_addrgen/$exit
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_word_addrgen/root_register_req
      -- CP-element group 175: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_word_addrgen/root_register_ack
      -- 
    ack_7400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx91_2830_delayed_6_0_2875_inst_ack_1, ack => convTransposeD_CP_6687_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	163 
    -- CP-element group 176: 	175 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/ptr_deref_2879_Split/$entry
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/ptr_deref_2879_Split/$exit
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/ptr_deref_2879_Split/split_req
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/ptr_deref_2879_Split/split_ack
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/word_access_start/$entry
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/word_access_start/word_0/$entry
      -- CP-element group 176: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/word_access_start/word_0/rr
      -- 
    rr_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(176), ack => ptr_deref_2879_store_0_req_0); -- 
    convTransposeD_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(163) & convTransposeD_CP_6687_elements(175) & convTransposeD_CP_6687_elements(178);
      gj_convTransposeD_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (5) 
      -- CP-element group 177: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/word_access_complete/word_0/cr
      -- CP-element group 177: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/word_access_complete/word_0/$entry
      -- CP-element group 177: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/word_access_complete/$entry
      -- CP-element group 177: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_update_start_
      -- CP-element group 177: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/$entry
      -- 
    cr_7449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(177), ack => ptr_deref_2879_store_0_req_1); -- 
    convTransposeD_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convTransposeD_CP_6687_elements(179);
      gj_convTransposeD_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	161 
    -- CP-element group 178: 	173 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (5) 
      -- CP-element group 178: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/word_access_start/$exit
      -- CP-element group 178: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/word_access_start/word_0/$exit
      -- CP-element group 178: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Sample/word_access_start/word_0/ra
      -- 
    ra_7439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2879_store_0_ack_0, ack => convTransposeD_CP_6687_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	209 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (5) 
      -- CP-element group 179: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/word_access_complete/word_0/ca
      -- CP-element group 179: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/word_access_complete/word_0/$exit
      -- CP-element group 179: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/word_access_complete/$exit
      -- CP-element group 179: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/ptr_deref_2879_Update/$exit
      -- 
    ca_7450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2879_store_0_ack_1, ack => convTransposeD_CP_6687_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	79 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_sample_start_
      -- 
    rr_7458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(180), ack => type_cast_2884_inst_req_0); -- 
    convTransposeD_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(79) & convTransposeD_CP_6687_elements(182);
      gj_convTransposeD_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	52 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	194 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_update_start_
      -- CP-element group 181: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Update/$entry
      -- 
    cr_7463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(181), ack => type_cast_2884_inst_req_1); -- 
    convTransposeD_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(183) & convTransposeD_CP_6687_elements(194);
      gj_convTransposeD_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	75 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Sample/ra
      -- 
    ra_7459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2884_inst_ack_0, ack => convTransposeD_CP_6687_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	192 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	74 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2884_Update/$exit
      -- 
    ca_7464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2884_inst_ack_1, ack => convTransposeD_CP_6687_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	49 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_sample_start_
      -- 
    rr_7472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(184), ack => type_cast_2888_inst_req_0); -- 
    convTransposeD_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(49) & convTransposeD_CP_6687_elements(186);
      gj_convTransposeD_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	52 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: 	194 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_update_start_
      -- 
    cr_7477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(185), ack => type_cast_2888_inst_req_1); -- 
    convTransposeD_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(187) & convTransposeD_CP_6687_elements(194);
      gj_convTransposeD_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_sample_completed_
      -- 
    ra_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2888_inst_ack_0, ack => convTransposeD_CP_6687_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	192 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	74 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2888_update_completed_
      -- 
    ca_7478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2888_inst_ack_1, ack => convTransposeD_CP_6687_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	79 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Sample/req
      -- CP-element group 188: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_sample_start_
      -- 
    req_7486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(188), ack => W_add106_2853_delayed_1_0_2902_inst_req_0); -- 
    convTransposeD_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(79) & convTransposeD_CP_6687_elements(190);
      gj_convTransposeD_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	52 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_update_start_
      -- CP-element group 189: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Update/req
      -- CP-element group 189: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Update/$entry
      -- 
    req_7491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(189), ack => W_add106_2853_delayed_1_0_2902_inst_req_1); -- 
    convTransposeD_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(191);
      gj_convTransposeD_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	75 
    -- CP-element group 190: 	188 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Sample/ack
      -- CP-element group 190: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_sample_completed_
      -- 
    ack_7487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add106_2853_delayed_1_0_2902_inst_ack_0, ack => convTransposeD_CP_6687_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	209 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	74 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Update/ack
      -- CP-element group 191: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2904_Update/$exit
      -- 
    ack_7492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add106_2853_delayed_1_0_2902_inst_ack_1, ack => convTransposeD_CP_6687_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	183 
    -- CP-element group 192: 	187 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_sample_start_
      -- 
    rr_7500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(192), ack => type_cast_2914_inst_req_0); -- 
    convTransposeD_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(183) & convTransposeD_CP_6687_elements(187) & convTransposeD_CP_6687_elements(194);
      gj_convTransposeD_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	52 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: 	202 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Update/cr
      -- CP-element group 193: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_update_start_
      -- 
    cr_7505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(193), ack => type_cast_2914_inst_req_1); -- 
    convTransposeD_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(195) & convTransposeD_CP_6687_elements(202);
      gj_convTransposeD_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	181 
    -- CP-element group 194: 	185 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_sample_completed_
      -- 
    ra_7501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_0, ack => convTransposeD_CP_6687_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	95 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2914_update_completed_
      -- 
    ca_7506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2914_inst_ack_1, ack => convTransposeD_CP_6687_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	100 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Sample/req
      -- CP-element group 196: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_sample_start_
      -- 
    req_7514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(196), ack => W_input_dim1x_x1_2870_delayed_2_0_2922_inst_req_0); -- 
    convTransposeD_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(100) & convTransposeD_CP_6687_elements(198);
      gj_convTransposeD_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	52 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	202 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Update/req
      -- CP-element group 197: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_update_start_
      -- 
    req_7519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(197), ack => W_input_dim1x_x1_2870_delayed_2_0_2922_inst_req_1); -- 
    convTransposeD_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(199) & convTransposeD_CP_6687_elements(202);
      gj_convTransposeD_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	96 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Sample/ack
      -- CP-element group 198: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_sample_completed_
      -- 
    ack_7515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_2870_delayed_2_0_2922_inst_ack_0, ack => convTransposeD_CP_6687_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	95 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Update/ack
      -- CP-element group 199: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2924_update_completed_
      -- 
    ack_7520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim1x_x1_2870_delayed_2_0_2922_inst_ack_1, ack => convTransposeD_CP_6687_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_sample_start_
      -- 
    rr_7528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(200), ack => type_cast_2937_inst_req_0); -- 
    convTransposeD_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(195) & convTransposeD_CP_6687_elements(199) & convTransposeD_CP_6687_elements(202);
      gj_convTransposeD_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	52 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Update/cr
      -- CP-element group 201: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_update_start_
      -- 
    cr_7533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(201), ack => type_cast_2937_inst_req_1); -- 
    convTransposeD_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(203);
      gj_convTransposeD_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	193 
    -- CP-element group 202: 	197 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_sample_completed_
      -- 
    ra_7529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2937_inst_ack_0, ack => convTransposeD_CP_6687_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	50 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	116 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Update/ca
      -- CP-element group 203: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/type_cast_2937_update_completed_
      -- 
    ca_7534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2937_inst_ack_1, ack => convTransposeD_CP_6687_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	121 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Sample/req
      -- CP-element group 204: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_sample_start_
      -- 
    req_7542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(204), ack => W_input_dim0x_x1_2884_delayed_3_0_2939_inst_req_0); -- 
    convTransposeD_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(121) & convTransposeD_CP_6687_elements(206);
      gj_convTransposeD_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	52 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Update/req
      -- CP-element group 205: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Update/$entry
      -- CP-element group 205: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_update_start_
      -- 
    req_7547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(205), ack => W_input_dim0x_x1_2884_delayed_3_0_2939_inst_req_1); -- 
    convTransposeD_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(207);
      gj_convTransposeD_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	117 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Sample/ack
      -- CP-element group 206: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_sample_completed_
      -- 
    ack_7543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_2884_delayed_3_0_2939_inst_ack_0, ack => convTransposeD_CP_6687_elements(206)); -- 
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	50 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	116 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Update/ack
      -- CP-element group 207: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/assign_stmt_2941_update_completed_
      -- 
    ack_7548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_dim0x_x1_2884_delayed_3_0_2939_inst_ack_1, ack => convTransposeD_CP_6687_elements(207)); -- 
    -- CP-element group 208:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	49 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	50 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convTransposeD_CP_6687_elements(208) is a control-delay.
    cp_element_208_delay: control_delay_element  generic map(name => " 208_delay", delay_value => 1)  port map(req => convTransposeD_CP_6687_elements(49), ack => convTransposeD_CP_6687_elements(208), clk => clk, reset =>reset);
    -- CP-element group 209:  join  transition  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	52 
    -- CP-element group 209: 	156 
    -- CP-element group 209: 	168 
    -- CP-element group 209: 	179 
    -- CP-element group 209: 	191 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	46 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_2618/do_while_stmt_2761/do_while_stmt_2761_loop_body/$exit
      -- 
    convTransposeD_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(52) & convTransposeD_CP_6687_elements(156) & convTransposeD_CP_6687_elements(168) & convTransposeD_CP_6687_elements(179) & convTransposeD_CP_6687_elements(191);
      gj_convTransposeD_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	45 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (2) 
      -- CP-element group 210: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_exit/ack
      -- CP-element group 210: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_exit/$exit
      -- 
    ack_7553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2761_branch_ack_0, ack => convTransposeD_CP_6687_elements(210)); -- 
    -- CP-element group 211:  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	45 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_taken/ack
      -- CP-element group 211: 	 branch_block_stmt_2618/do_while_stmt_2761/loop_taken/$exit
      -- 
    ack_7557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2761_branch_ack_1, ack => convTransposeD_CP_6687_elements(211)); -- 
    -- CP-element group 212:  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	43 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	1 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_2618/do_while_stmt_2761/$exit
      -- 
    convTransposeD_CP_6687_elements(212) <= convTransposeD_CP_6687_elements(43);
    -- CP-element group 213:  merge  transition  place  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	1 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (15) 
      -- CP-element group 213: 	 branch_block_stmt_2618/merge_stmt_2975__exit__
      -- CP-element group 213: 	 branch_block_stmt_2618/assign_stmt_2980__entry__
      -- CP-element group 213: 	 branch_block_stmt_2618/assign_stmt_2980/$entry
      -- CP-element group 213: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_sample_start_
      -- CP-element group 213: 	 branch_block_stmt_2618/merge_stmt_2975_PhiReqMerge
      -- CP-element group 213: 	 branch_block_stmt_2618/whilex_xbody_whilex_xend
      -- CP-element group 213: 	 branch_block_stmt_2618/if_stmt_2971_if_link/if_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_2618/if_stmt_2971_if_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Sample/req
      -- CP-element group 213: 	 branch_block_stmt_2618/merge_stmt_2975_PhiAck/dummy
      -- CP-element group 213: 	 branch_block_stmt_2618/merge_stmt_2975_PhiAck/$exit
      -- CP-element group 213: 	 branch_block_stmt_2618/merge_stmt_2975_PhiAck/$entry
      -- CP-element group 213: 	 branch_block_stmt_2618/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 213: 	 branch_block_stmt_2618/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Sample/$entry
      -- 
    if_choice_transition_7571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2971_branch_ack_1, ack => convTransposeD_CP_6687_elements(213)); -- 
    req_7587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(213), ack => WPIPE_Block3_done_2977_inst_req_0); -- 
    -- CP-element group 214:  merge  transition  place  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	1 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (5) 
      -- CP-element group 214: 	 branch_block_stmt_2618/if_stmt_2971__exit__
      -- CP-element group 214: 	 branch_block_stmt_2618/merge_stmt_2975__entry__
      -- CP-element group 214: 	 branch_block_stmt_2618/if_stmt_2971_else_link/else_choice_transition
      -- CP-element group 214: 	 branch_block_stmt_2618/if_stmt_2971_else_link/$exit
      -- CP-element group 214: 	 branch_block_stmt_2618/merge_stmt_2975_dead_link/$entry
      -- 
    else_choice_transition_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2971_branch_ack_0, ack => convTransposeD_CP_6687_elements(214)); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Update/req
      -- CP-element group 215: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_update_start_
      -- CP-element group 215: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_sample_completed_
      -- 
    ack_7588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2977_inst_ack_0, ack => convTransposeD_CP_6687_elements(215)); -- 
    req_7592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(215), ack => WPIPE_Block3_done_2977_inst_req_1); -- 
    -- CP-element group 216:  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (16) 
      -- CP-element group 216: 	 branch_block_stmt_2618/branch_block_stmt_2618__exit__
      -- CP-element group 216: 	 $exit
      -- CP-element group 216: 	 branch_block_stmt_2618/$exit
      -- CP-element group 216: 	 branch_block_stmt_2618/assign_stmt_2980__exit__
      -- CP-element group 216: 	 branch_block_stmt_2618/return__
      -- CP-element group 216: 	 branch_block_stmt_2618/merge_stmt_2982__exit__
      -- CP-element group 216: 	 branch_block_stmt_2618/assign_stmt_2980/$exit
      -- CP-element group 216: 	 branch_block_stmt_2618/merge_stmt_2982_PhiReqMerge
      -- CP-element group 216: 	 branch_block_stmt_2618/merge_stmt_2982_PhiAck/dummy
      -- CP-element group 216: 	 branch_block_stmt_2618/merge_stmt_2982_PhiAck/$exit
      -- CP-element group 216: 	 branch_block_stmt_2618/merge_stmt_2982_PhiAck/$entry
      -- CP-element group 216: 	 branch_block_stmt_2618/return___PhiReq/$exit
      -- CP-element group 216: 	 branch_block_stmt_2618/return___PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Update/ack
      -- CP-element group 216: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_2618/assign_stmt_2980/WPIPE_Block3_done_2977_update_completed_
      -- 
    ack_7593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2977_inst_ack_1, ack => convTransposeD_CP_6687_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	41 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (2) 
      -- CP-element group 217: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Sample/$exit
      -- 
    ra_7613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2759_inst_ack_0, ack => convTransposeD_CP_6687_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	41 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/ca
      -- CP-element group 218: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/Update/$exit
      -- 
    ca_7618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2759_inst_ack_1, ack => convTransposeD_CP_6687_elements(218)); -- 
    -- CP-element group 219:  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (8) 
      -- CP-element group 219: 	 branch_block_stmt_2618/merge_stmt_2740_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_req
      -- CP-element group 219: 	 branch_block_stmt_2618/merge_stmt_2740_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/SplitProtocol/$exit
      -- CP-element group 219: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/type_cast_2759/$exit
      -- CP-element group 219: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/phi_stmt_2756_sources/$exit
      -- CP-element group 219: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/phi_stmt_2756/$exit
      -- CP-element group 219: 	 branch_block_stmt_2618/entry_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2756_req_7619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2756_req_7619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6687_elements(219), ack => phi_stmt_2756_req_0); -- 
    convTransposeD_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6687_elements(217) & convTransposeD_CP_6687_elements(218);
      gj_convTransposeD_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6687_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	42 
    -- CP-element group 220:  members (4) 
      -- CP-element group 220: 	 branch_block_stmt_2618/do_while_stmt_2761__entry__
      -- CP-element group 220: 	 branch_block_stmt_2618/merge_stmt_2740__exit__
      -- CP-element group 220: 	 branch_block_stmt_2618/merge_stmt_2740_PhiAck/$exit
      -- CP-element group 220: 	 branch_block_stmt_2618/merge_stmt_2740_PhiAck/phi_stmt_2756_ack
      -- 
    phi_stmt_2756_ack_7624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2756_ack_0, ack => convTransposeD_CP_6687_elements(220)); -- 
    convTransposeD_do_while_stmt_2761_terminator_7558: loop_terminator -- 
      generic map (name => " convTransposeD_do_while_stmt_2761_terminator_7558", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convTransposeD_CP_6687_elements(46),loop_continue => convTransposeD_CP_6687_elements(211),loop_terminate => convTransposeD_CP_6687_elements(210),loop_back => convTransposeD_CP_6687_elements(44),loop_exit => convTransposeD_CP_6687_elements(43),clk => clk, reset => reset); -- 
    phi_stmt_2763_phi_seq_7046_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeD_CP_6687_elements(59);
      convTransposeD_CP_6687_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeD_CP_6687_elements(68);
      convTransposeD_CP_6687_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeD_CP_6687_elements(69);
      convTransposeD_CP_6687_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeD_CP_6687_elements(61);
      convTransposeD_CP_6687_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeD_CP_6687_elements(70);
      convTransposeD_CP_6687_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeD_CP_6687_elements(72);
      convTransposeD_CP_6687_elements(62) <= phi_mux_reqs(1);
      phi_stmt_2763_phi_seq_7046 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2763_phi_seq_7046") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeD_CP_6687_elements(51), 
          phi_sample_ack => convTransposeD_CP_6687_elements(57), 
          phi_update_req => convTransposeD_CP_6687_elements(53), 
          phi_update_ack => convTransposeD_CP_6687_elements(58), 
          phi_mux_ack => convTransposeD_CP_6687_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2768_phi_seq_7090_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeD_CP_6687_elements(80);
      convTransposeD_CP_6687_elements(85)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeD_CP_6687_elements(89);
      convTransposeD_CP_6687_elements(86)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeD_CP_6687_elements(90);
      convTransposeD_CP_6687_elements(81) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeD_CP_6687_elements(82);
      convTransposeD_CP_6687_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeD_CP_6687_elements(91);
      convTransposeD_CP_6687_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeD_CP_6687_elements(93);
      convTransposeD_CP_6687_elements(83) <= phi_mux_reqs(1);
      phi_stmt_2768_phi_seq_7090 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2768_phi_seq_7090") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeD_CP_6687_elements(76), 
          phi_sample_ack => convTransposeD_CP_6687_elements(77), 
          phi_update_req => convTransposeD_CP_6687_elements(78), 
          phi_update_ack => convTransposeD_CP_6687_elements(79), 
          phi_mux_ack => convTransposeD_CP_6687_elements(84), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2773_phi_seq_7134_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeD_CP_6687_elements(101);
      convTransposeD_CP_6687_elements(106)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeD_CP_6687_elements(110);
      convTransposeD_CP_6687_elements(107)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeD_CP_6687_elements(111);
      convTransposeD_CP_6687_elements(102) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeD_CP_6687_elements(103);
      convTransposeD_CP_6687_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeD_CP_6687_elements(112);
      convTransposeD_CP_6687_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeD_CP_6687_elements(114);
      convTransposeD_CP_6687_elements(104) <= phi_mux_reqs(1);
      phi_stmt_2773_phi_seq_7134 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2773_phi_seq_7134") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeD_CP_6687_elements(97), 
          phi_sample_ack => convTransposeD_CP_6687_elements(98), 
          phi_update_req => convTransposeD_CP_6687_elements(99), 
          phi_update_ack => convTransposeD_CP_6687_elements(100), 
          phi_mux_ack => convTransposeD_CP_6687_elements(105), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2778_phi_seq_7188_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convTransposeD_CP_6687_elements(122);
      convTransposeD_CP_6687_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convTransposeD_CP_6687_elements(131);
      convTransposeD_CP_6687_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= convTransposeD_CP_6687_elements(132);
      convTransposeD_CP_6687_elements(123) <= phi_mux_reqs(0);
      triggers(1)  <= convTransposeD_CP_6687_elements(124);
      convTransposeD_CP_6687_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convTransposeD_CP_6687_elements(135);
      convTransposeD_CP_6687_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= convTransposeD_CP_6687_elements(136);
      convTransposeD_CP_6687_elements(125) <= phi_mux_reqs(1);
      phi_stmt_2778_phi_seq_7188 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2778_phi_seq_7188") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convTransposeD_CP_6687_elements(118), 
          phi_sample_ack => convTransposeD_CP_6687_elements(119), 
          phi_update_req => convTransposeD_CP_6687_elements(120), 
          phi_update_ack => convTransposeD_CP_6687_elements(121), 
          phi_mux_ack => convTransposeD_CP_6687_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6998_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convTransposeD_CP_6687_elements(47);
        preds(1)  <= convTransposeD_CP_6687_elements(48);
        entry_tmerge_6998 : transition_merge -- 
          generic map(name => " entry_tmerge_6998")
          port map (preds => preds, symbol_out => convTransposeD_CP_6687_elements(49));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_2970_wire : std_logic_vector(0 downto 0);
    signal R_idxprom90_2871_resized : std_logic_vector(13 downto 0);
    signal R_idxprom90_2871_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2848_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2848_scaled : std_logic_vector(13 downto 0);
    signal add106_2853_delayed_1_0_2904 : std_logic_vector(15 downto 0);
    signal add106_2901 : std_logic_vector(15 downto 0);
    signal add32_2697 : std_logic_vector(15 downto 0);
    signal add50_2703 : std_logic_vector(15 downto 0);
    signal add63_2714 : std_logic_vector(15 downto 0);
    signal add82_2830 : std_logic_vector(63 downto 0);
    signal add84_2840 : std_logic_vector(63 downto 0);
    signal add_2670 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2788 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2849_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2849_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2849_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2849_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2849_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2849_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2872_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2872_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2872_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2872_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2872_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2872_root_address : std_logic_vector(13 downto 0);
    signal arrayidx86_2851 : std_logic_vector(31 downto 0);
    signal arrayidx91_2830_delayed_6_0_2877 : std_logic_vector(31 downto 0);
    signal arrayidx91_2874 : std_logic_vector(31 downto 0);
    signal call11_2639 : std_logic_vector(15 downto 0);
    signal call13_2642 : std_logic_vector(15 downto 0);
    signal call14_2645 : std_logic_vector(15 downto 0);
    signal call15_2648 : std_logic_vector(15 downto 0);
    signal call16_2661 : std_logic_vector(15 downto 0);
    signal call18_2673 : std_logic_vector(15 downto 0);
    signal call1_2624 : std_logic_vector(15 downto 0);
    signal call20_2676 : std_logic_vector(15 downto 0);
    signal call22_2679 : std_logic_vector(15 downto 0);
    signal call3_2627 : std_logic_vector(15 downto 0);
    signal call5_2630 : std_logic_vector(15 downto 0);
    signal call7_2633 : std_logic_vector(15 downto 0);
    signal call9_2636 : std_logic_vector(15 downto 0);
    signal call_2621 : std_logic_vector(15 downto 0);
    signal cmp114_2934 : std_logic_vector(0 downto 0);
    signal cmp125_2958 : std_logic_vector(0 downto 0);
    signal cmp_2895 : std_logic_vector(0 downto 0);
    signal conv100_2885 : std_logic_vector(31 downto 0);
    signal conv102_2738 : std_logic_vector(31 downto 0);
    signal conv17_2665 : std_logic_vector(31 downto 0);
    signal conv70_2812 : std_logic_vector(63 downto 0);
    signal conv73_2723 : std_logic_vector(63 downto 0);
    signal conv75_2816 : std_logic_vector(63 downto 0);
    signal conv78_2727 : std_logic_vector(63 downto 0);
    signal conv80_2820 : std_logic_vector(63 downto 0);
    signal conv_2652 : std_logic_vector(31 downto 0);
    signal iNsTr_18_2915 : std_logic_vector(15 downto 0);
    signal idxprom90_2867 : std_logic_vector(63 downto 0);
    signal idxprom_2844 : std_logic_vector(63 downto 0);
    signal inc118_2938 : std_logic_vector(15 downto 0);
    signal inc118x_xinput_dim0x_x1_2946 : std_logic_vector(15 downto 0);
    signal inc_2921 : std_logic_vector(15 downto 0);
    signal indvar_2763 : std_logic_vector(31 downto 0);
    signal indvar_at_entry_2741 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2964 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1_2778 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_2884_delayed_3_0_2941 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_2756 : std_logic_vector(15 downto 0);
    signal input_dim0x_x1_at_entry_2756_2782_buffered : std_logic_vector(15 downto 0);
    signal input_dim1x_x0_2929 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2773 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2870_delayed_2_0_2924 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_at_entry_2751 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2953 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0_2911 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2768 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_at_entry_2746 : std_logic_vector(15 downto 0);
    signal mul59_2803 : std_logic_vector(15 downto 0);
    signal mul81_2825 : std_logic_vector(63 downto 0);
    signal mul83_2835 : std_logic_vector(63 downto 0);
    signal mul_2793 : std_logic_vector(15 downto 0);
    signal ptr_deref_2854_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2854_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2854_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2854_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2854_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2879_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2879_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2879_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2879_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2879_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2879_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2658 : std_logic_vector(31 downto 0);
    signal shr138_2686 : std_logic_vector(15 downto 0);
    signal shr31139_2692 : std_logic_vector(15 downto 0);
    signal shr89_2861 : std_logic_vector(63 downto 0);
    signal sub53_2798 : std_logic_vector(15 downto 0);
    signal sub66_2719 : std_logic_vector(15 downto 0);
    signal sub67_2808 : std_logic_vector(15 downto 0);
    signal sub96_2733 : std_logic_vector(15 downto 0);
    signal sub_2708 : std_logic_vector(15 downto 0);
    signal tmp87_2855 : std_logic_vector(63 downto 0);
    signal type_cast_2656_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2684_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2690_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2701_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2712_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2731_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2736_wire : std_logic_vector(31 downto 0);
    signal type_cast_2759_wire : std_logic_vector(15 downto 0);
    signal type_cast_2766_wire : std_logic_vector(31 downto 0);
    signal type_cast_2771_wire : std_logic_vector(15 downto 0);
    signal type_cast_2776_wire : std_logic_vector(15 downto 0);
    signal type_cast_2781_wire : std_logic_vector(15 downto 0);
    signal type_cast_2842_2842_delayed_2_0_2889 : std_logic_vector(31 downto 0);
    signal type_cast_2859_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2865_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2892_wire : std_logic_vector(31 downto 0);
    signal type_cast_2899_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2909_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2919_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2950_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2979_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_whilex_xend_taken_2967 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_2849_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2849_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2849_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2849_resized_base_address <= "00000000000000";
    array_obj_ref_2872_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2872_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2872_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2872_resized_base_address <= "00000000000000";
    indvar_at_entry_2741 <= "00000000000000000000000000000000";
    input_dim1x_x1_at_entry_2751 <= "0000000000000000";
    input_dim2x_x1_at_entry_2746 <= "0000000000000000";
    ptr_deref_2854_word_offset_0 <= "00000000000000";
    ptr_deref_2879_word_offset_0 <= "00000000000000";
    type_cast_2656_wire_constant <= "00000000000000000000000000010000";
    type_cast_2684_wire_constant <= "0000000000000010";
    type_cast_2690_wire_constant <= "0000000000000001";
    type_cast_2701_wire_constant <= "1111111111111111";
    type_cast_2712_wire_constant <= "1111111111111111";
    type_cast_2731_wire_constant <= "1111111111111100";
    type_cast_2859_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2865_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2899_wire_constant <= "0000000000000100";
    type_cast_2909_wire_constant <= "0000000000000000";
    type_cast_2919_wire_constant <= "0000000000000001";
    type_cast_2950_wire_constant <= "0000000000000000";
    type_cast_2962_wire_constant <= "00000000000000000000000000000001";
    type_cast_2979_wire_constant <= "0000000000000001";
    phi_stmt_2756: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2759_wire;
      req(0) <= phi_stmt_2756_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2756",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2756_ack_0,
          idata => idata,
          odata => input_dim0x_x1_at_entry_2756,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2756
    phi_stmt_2763: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2766_wire & indvar_at_entry_2741;
      req <= phi_stmt_2763_req_0 & phi_stmt_2763_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2763",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2763_ack_0,
          idata => idata,
          odata => indvar_2763,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2763
    phi_stmt_2768: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2771_wire & input_dim2x_x1_at_entry_2746;
      req <= phi_stmt_2768_req_0 & phi_stmt_2768_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2768",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2768_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2768,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2768
    phi_stmt_2773: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2776_wire & input_dim1x_x1_at_entry_2751;
      req <= phi_stmt_2773_req_0 & phi_stmt_2773_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2773",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2773_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2773,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2773
    phi_stmt_2778: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2781_wire & input_dim0x_x1_at_entry_2756_2782_buffered;
      req <= phi_stmt_2778_req_0 & phi_stmt_2778_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2778",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2778_ack_0,
          idata => idata,
          odata => input_dim0x_x1_2778,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2778
    -- flow-through select operator MUX_2910_inst
    input_dim2x_x0_2911 <= add106_2853_delayed_1_0_2904 when (cmp_2895(0) /=  '0') else type_cast_2909_wire_constant;
    -- flow-through select operator MUX_2952_inst
    input_dim1x_x2_2953 <= type_cast_2950_wire_constant when (cmp114_2934(0) /=  '0') else input_dim1x_x0_2929;
    W_add106_2853_delayed_1_0_2902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add106_2853_delayed_1_0_2902_inst_req_0;
      W_add106_2853_delayed_1_0_2902_inst_ack_0<= wack(0);
      rreq(0) <= W_add106_2853_delayed_1_0_2902_inst_req_1;
      W_add106_2853_delayed_1_0_2902_inst_ack_1<= rack(0);
      W_add106_2853_delayed_1_0_2902_inst : InterlockBuffer generic map ( -- 
        name => "W_add106_2853_delayed_1_0_2902_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add106_2901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add106_2853_delayed_1_0_2904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx91_2830_delayed_6_0_2875_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx91_2830_delayed_6_0_2875_inst_req_0;
      W_arrayidx91_2830_delayed_6_0_2875_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx91_2830_delayed_6_0_2875_inst_req_1;
      W_arrayidx91_2830_delayed_6_0_2875_inst_ack_1<= rack(0);
      W_arrayidx91_2830_delayed_6_0_2875_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx91_2830_delayed_6_0_2875_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx91_2874,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx91_2830_delayed_6_0_2877,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim0x_x1_2884_delayed_3_0_2939_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim0x_x1_2884_delayed_3_0_2939_inst_req_0;
      W_input_dim0x_x1_2884_delayed_3_0_2939_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim0x_x1_2884_delayed_3_0_2939_inst_req_1;
      W_input_dim0x_x1_2884_delayed_3_0_2939_inst_ack_1<= rack(0);
      W_input_dim0x_x1_2884_delayed_3_0_2939_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim0x_x1_2884_delayed_3_0_2939_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_2778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_2884_delayed_3_0_2941,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_dim1x_x1_2870_delayed_2_0_2922_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_dim1x_x1_2870_delayed_2_0_2922_inst_req_0;
      W_input_dim1x_x1_2870_delayed_2_0_2922_inst_ack_0<= wack(0);
      rreq(0) <= W_input_dim1x_x1_2870_delayed_2_0_2922_inst_req_1;
      W_input_dim1x_x1_2870_delayed_2_0_2922_inst_ack_1<= rack(0);
      W_input_dim1x_x1_2870_delayed_2_0_2922_inst : InterlockBuffer generic map ( -- 
        name => "W_input_dim1x_x1_2870_delayed_2_0_2922_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2773,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim1x_x1_2870_delayed_2_0_2924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_2965_inst
    process(cmp125_2958) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp125_2958(0 downto 0);
      whilex_xbody_whilex_xend_taken_2967 <= tmp_var; -- 
    end process;
    addr_of_2850_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2850_final_reg_req_0;
      addr_of_2850_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2850_final_reg_req_1;
      addr_of_2850_final_reg_ack_1<= rack(0);
      addr_of_2850_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2850_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2849_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx86_2851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2873_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2873_final_reg_req_0;
      addr_of_2873_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2873_final_reg_req_1;
      addr_of_2873_final_reg_ack_1<= rack(0);
      addr_of_2873_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2873_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2872_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx91_2874,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    input_dim0x_x1_at_entry_2756_2782_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= input_dim0x_x1_at_entry_2756_2782_buf_req_0;
      input_dim0x_x1_at_entry_2756_2782_buf_ack_0<= wack(0);
      rreq(0) <= input_dim0x_x1_at_entry_2756_2782_buf_req_1;
      input_dim0x_x1_at_entry_2756_2782_buf_ack_1<= rack(0);
      input_dim0x_x1_at_entry_2756_2782_buf : InterlockBuffer generic map ( -- 
        name => "input_dim0x_x1_at_entry_2756_2782_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1_at_entry_2756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_dim0x_x1_at_entry_2756_2782_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2651_inst_req_0;
      type_cast_2651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2651_inst_req_1;
      type_cast_2651_inst_ack_1<= rack(0);
      type_cast_2651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2664_inst_req_0;
      type_cast_2664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2664_inst_req_1;
      type_cast_2664_inst_ack_1<= rack(0);
      type_cast_2664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2722_inst_req_0;
      type_cast_2722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2722_inst_req_1;
      type_cast_2722_inst_ack_1<= rack(0);
      type_cast_2722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2679,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2726_inst_req_0;
      type_cast_2726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2726_inst_req_1;
      type_cast_2726_inst_ack_1<= rack(0);
      type_cast_2726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2737_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2737_inst_req_0;
      type_cast_2737_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2737_inst_req_1;
      type_cast_2737_inst_ack_1<= rack(0);
      type_cast_2737_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2737_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2736_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_2738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2759_inst_req_0;
      type_cast_2759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2759_inst_req_1;
      type_cast_2759_inst_ack_1<= rack(0);
      type_cast_2759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2759_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2697,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2759_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2766_inst_req_0;
      type_cast_2766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2766_inst_req_1;
      type_cast_2766_inst_ack_1<= rack(0);
      type_cast_2766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2766_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2964,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2766_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2771_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2771_inst_req_0;
      type_cast_2771_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2771_inst_req_1;
      type_cast_2771_inst_ack_1<= rack(0);
      type_cast_2771_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2771_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0_2911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2771_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2776_inst_req_0;
      type_cast_2776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2776_inst_req_1;
      type_cast_2776_inst_ack_1<= rack(0);
      type_cast_2776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2776_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2953,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2776_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2781_inst_req_0;
      type_cast_2781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2781_inst_req_1;
      type_cast_2781_inst_ack_1<= rack(0);
      type_cast_2781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2781_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc118x_xinput_dim0x_x1_2946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2781_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2811_inst_req_0;
      type_cast_2811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2811_inst_req_1;
      type_cast_2811_inst_ack_1<= rack(0);
      type_cast_2811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2812,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2815_inst_req_0;
      type_cast_2815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2815_inst_req_1;
      type_cast_2815_inst_ack_1<= rack(0);
      type_cast_2815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2819_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2819_inst_req_0;
      type_cast_2819_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2819_inst_req_1;
      type_cast_2819_inst_ack_1<= rack(0);
      type_cast_2819_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2819_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2820,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2843_inst_req_0;
      type_cast_2843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2843_inst_req_1;
      type_cast_2843_inst_ack_1<= rack(0);
      type_cast_2843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_src_0x_x0_2788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2884_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2884_inst_req_0;
      type_cast_2884_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2884_inst_req_1;
      type_cast_2884_inst_ack_1<= rack(0);
      type_cast_2884_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2884_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_2885,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2888_inst_req_0;
      type_cast_2888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2888_inst_req_1;
      type_cast_2888_inst_ack_1<= rack(0);
      type_cast_2888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2888_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv102_2738,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2842_2842_delayed_2_0_2889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2892_inst
    process(conv100_2885) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv100_2885(31 downto 0);
      type_cast_2892_wire <= tmp_var; -- 
    end process;
    type_cast_2914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2914_inst_req_0;
      type_cast_2914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2914_inst_req_1;
      type_cast_2914_inst_ack_1<= rack(0);
      type_cast_2914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2914_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_2895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_18_2915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2937_inst_req_0;
      type_cast_2937_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2937_inst_req_1;
      type_cast_2937_inst_ack_1<= rack(0);
      type_cast_2937_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2937_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp114_2934,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc118_2938,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2849_index_1_rename
    process(R_idxprom_2848_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2848_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2848_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2849_index_1_resize
    process(idxprom_2844) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2844;
      ov := iv(13 downto 0);
      R_idxprom_2848_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2849_root_address_inst
    process(array_obj_ref_2849_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2849_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2849_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2872_index_1_rename
    process(R_idxprom90_2871_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom90_2871_resized;
      ov(13 downto 0) := iv;
      R_idxprom90_2871_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2872_index_1_resize
    process(idxprom90_2867) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom90_2867;
      ov := iv(13 downto 0);
      R_idxprom90_2871_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2872_root_address_inst
    process(array_obj_ref_2872_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2872_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2872_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2854_addr_0
    process(ptr_deref_2854_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2854_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2854_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2854_base_resize
    process(arrayidx86_2851) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx86_2851;
      ov := iv(13 downto 0);
      ptr_deref_2854_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2854_gather_scatter
    process(ptr_deref_2854_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2854_data_0;
      ov(63 downto 0) := iv;
      tmp87_2855 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2854_root_address_inst
    process(ptr_deref_2854_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2854_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2854_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2879_addr_0
    process(ptr_deref_2879_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2879_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2879_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2879_base_resize
    process(arrayidx91_2830_delayed_6_0_2877) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx91_2830_delayed_6_0_2877;
      ov := iv(13 downto 0);
      ptr_deref_2879_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2879_gather_scatter
    process(tmp87_2855) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp87_2855;
      ov(63 downto 0) := iv;
      ptr_deref_2879_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2879_root_address_inst
    process(ptr_deref_2879_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2879_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2879_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_2761_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2970_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2761_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2761_branch_req_0,
          ack0 => do_while_stmt_2761_branch_ack_0,
          ack1 => do_while_stmt_2761_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2971_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_2967;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2971_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2971_branch_req_0,
          ack0 => if_stmt_2971_branch_ack_0,
          ack1 => if_stmt_2971_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2696_inst
    process(shr138_2686, shr31139_2692) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr138_2686, shr31139_2692, tmp_var);
      add32_2697 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2702_inst
    process(call7_2633) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2633, type_cast_2701_wire_constant, tmp_var);
      add50_2703 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2713_inst
    process(call9_2636) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2636, type_cast_2712_wire_constant, tmp_var);
      add63_2714 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2732_inst
    process(call3_2627) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call3_2627, type_cast_2731_wire_constant, tmp_var);
      sub96_2733 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2797_inst
    process(sub_2708, mul_2793) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2708, mul_2793, tmp_var);
      sub53_2798 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2807_inst
    process(sub66_2719, mul59_2803) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2719, mul59_2803, tmp_var);
      sub67_2808 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2900_inst
    process(input_dim2x_x1_2768) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2768, type_cast_2899_wire_constant, tmp_var);
      add106_2901 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2928_inst
    process(inc_2921, input_dim1x_x1_2870_delayed_2_0_2924) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc_2921, input_dim1x_x1_2870_delayed_2_0_2924, tmp_var);
      input_dim1x_x0_2929 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2945_inst
    process(inc118_2938, input_dim0x_x1_2884_delayed_3_0_2941) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc118_2938, input_dim0x_x1_2884_delayed_3_0_2941, tmp_var);
      inc118x_xinput_dim0x_x1_2946 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2787_inst
    process(add_2670, indvar_2763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2670, indvar_2763, tmp_var);
      add_src_0x_x0_2788 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2963_inst
    process(indvar_2763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2763, type_cast_2962_wire_constant, tmp_var);
      indvarx_xnext_2964 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2829_inst
    process(mul81_2825, conv75_2816) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2825, conv75_2816, tmp_var);
      add82_2830 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2839_inst
    process(mul83_2835, conv70_2812) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2835, conv70_2812, tmp_var);
      add84_2840 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2866_inst
    process(shr89_2861) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr89_2861, type_cast_2865_wire_constant, tmp_var);
      idxprom90_2867 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2933_inst
    process(input_dim1x_x0_2929, call1_2624) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1x_x0_2929, call1_2624, tmp_var);
      cmp114_2934 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2957_inst
    process(inc118x_xinput_dim0x_x1_2946, call_2621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc118x_xinput_dim0x_x1_2946, call_2621, tmp_var);
      cmp125_2958 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2685_inst
    process(call_2621) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2621, type_cast_2684_wire_constant, tmp_var);
      shr138_2686 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2691_inst
    process(call_2621) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2621, type_cast_2690_wire_constant, tmp_var);
      shr31139_2692 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2860_inst
    process(add84_2840) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2840, type_cast_2859_wire_constant, tmp_var);
      shr89_2861 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2792_inst
    process(input_dim0x_x1_2778, call13_2642) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x1_2778, call13_2642, tmp_var);
      mul_2793 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2802_inst
    process(input_dim1x_x1_2773, call13_2642) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2773, call13_2642, tmp_var);
      mul59_2803 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2824_inst
    process(conv80_2820, conv78_2727) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2820, conv78_2727, tmp_var);
      mul81_2825 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2834_inst
    process(add82_2830, conv73_2723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2830, conv73_2723, tmp_var);
      mul83_2835 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2970_inst
    process(cmp125_2958) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp125_2958, tmp_var);
      NOT_u1_u1_2970_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u32_u32_2669_inst
    process(shl_2658, conv17_2665) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2658, conv17_2665, tmp_var);
      add_2670 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2657_inst
    process(conv_2652) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2652, type_cast_2656_wire_constant, tmp_var);
      shl_2658 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2894_inst
    process(type_cast_2892_wire, type_cast_2842_2842_delayed_2_0_2889) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2892_wire, type_cast_2842_2842_delayed_2_0_2889, tmp_var);
      cmp_2895 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2707_inst
    process(add50_2703, call14_2645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2703, call14_2645, tmp_var);
      sub_2708 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2718_inst
    process(add63_2714, call14_2645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2714, call14_2645, tmp_var);
      sub66_2719 <= tmp_var; --
    end process;
    -- binary operator XOR_u16_u16_2920_inst
    process(iNsTr_18_2915) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntXor_proc(iNsTr_18_2915, type_cast_2919_wire_constant, tmp_var);
      inc_2921 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2849_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2848_scaled;
      array_obj_ref_2849_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2849_index_offset_req_0;
      array_obj_ref_2849_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2849_index_offset_req_1;
      array_obj_ref_2849_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2872_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom90_2871_scaled;
      array_obj_ref_2872_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2872_index_offset_req_0;
      array_obj_ref_2872_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2872_index_offset_req_1;
      array_obj_ref_2872_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- unary operator type_cast_2736_inst
    process(sub96_2733) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", sub96_2733, tmp_var);
      type_cast_2736_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_2854_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2854_load_0_req_0;
      ptr_deref_2854_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2854_load_0_req_1;
      ptr_deref_2854_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2854_word_address_0;
      ptr_deref_2854_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2879_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 15);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2879_store_0_req_0;
      ptr_deref_2879_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2879_store_0_req_1;
      ptr_deref_2879_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2879_word_address_0;
      data_in <= ptr_deref_2879_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2620_inst RPIPE_Block3_start_2626_inst RPIPE_Block3_start_2641_inst RPIPE_Block3_start_2647_inst RPIPE_Block3_start_2644_inst RPIPE_Block3_start_2623_inst RPIPE_Block3_start_2638_inst RPIPE_Block3_start_2678_inst RPIPE_Block3_start_2672_inst RPIPE_Block3_start_2660_inst RPIPE_Block3_start_2635_inst RPIPE_Block3_start_2675_inst RPIPE_Block3_start_2632_inst RPIPE_Block3_start_2629_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2620_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2626_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2641_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2647_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2644_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2623_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2638_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2678_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2672_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2660_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2635_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2675_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2632_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2629_inst_req_0;
      RPIPE_Block3_start_2620_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2626_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2641_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2647_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2644_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2623_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2638_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2678_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2672_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2660_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2635_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2675_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2632_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2629_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2620_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2626_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2641_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2647_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2644_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2623_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2638_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2678_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2672_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2660_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2635_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2675_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2632_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2629_inst_req_1;
      RPIPE_Block3_start_2620_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2626_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2641_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2647_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2644_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2623_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2638_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2678_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2672_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2660_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2635_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2675_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2632_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2629_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2621 <= data_out(223 downto 208);
      call3_2627 <= data_out(207 downto 192);
      call13_2642 <= data_out(191 downto 176);
      call15_2648 <= data_out(175 downto 160);
      call14_2645 <= data_out(159 downto 144);
      call1_2624 <= data_out(143 downto 128);
      call11_2639 <= data_out(127 downto 112);
      call22_2679 <= data_out(111 downto 96);
      call18_2673 <= data_out(95 downto 80);
      call16_2661 <= data_out(79 downto 64);
      call9_2636 <= data_out(63 downto 48);
      call20_2676 <= data_out(47 downto 32);
      call7_2633 <= data_out(31 downto 16);
      call5_2630 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2977_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2977_inst_req_0;
      WPIPE_Block3_done_2977_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2977_inst_req_1;
      WPIPE_Block3_done_2977_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2979_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_resp_34_inst_req_0 : boolean;
  signal RPIPE_timer_resp_34_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_34_inst_req_1 : boolean;
  signal RPIPE_timer_resp_34_inst_ack_1 : boolean;
  signal WPIPE_timer_req_29_inst_req_0 : boolean;
  signal WPIPE_timer_req_29_inst_ack_0 : boolean;
  signal WPIPE_timer_req_29_inst_req_1 : boolean;
  signal WPIPE_timer_req_29_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_sample_start_
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/req
      -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_29_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_34_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_update_start_
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/ack
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/$entry
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_29_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_29_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_29_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_sample_completed_
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_update_start_
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/ra
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/$entry
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_34_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_34_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_update_completed_
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/$exit
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_34_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_32_to_assign_stmt_35/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(4) & timer_CP_0_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_31_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_31_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_34_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_34_inst_req_0;
      RPIPE_timer_resp_34_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_34_inst_req_1;
      RPIPE_timer_resp_34_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_29_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_29_inst_req_0;
      WPIPE_timer_req_29_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_29_inst_req_1;
      WPIPE_timer_req_29_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_31_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_7671_start: Boolean;
  signal timerDaemon_CP_7671_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_req_3004_inst_ack_1 : boolean;
  signal do_while_stmt_2995_branch_req_0 : boolean;
  signal WPIPE_timer_resp_3012_inst_req_1 : boolean;
  signal WPIPE_timer_resp_3012_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_3012_inst_req_0 : boolean;
  signal nCOUNTER_3010_3001_buf_req_1 : boolean;
  signal nCOUNTER_3010_3001_buf_ack_1 : boolean;
  signal phi_stmt_2997_req_1 : boolean;
  signal phi_stmt_2997_req_0 : boolean;
  signal RPIPE_timer_req_3004_inst_req_0 : boolean;
  signal do_while_stmt_2995_branch_ack_0 : boolean;
  signal WPIPE_timer_resp_3012_inst_ack_0 : boolean;
  signal nCOUNTER_3010_3001_buf_req_0 : boolean;
  signal nCOUNTER_3010_3001_buf_ack_0 : boolean;
  signal RPIPE_timer_req_3004_inst_req_1 : boolean;
  signal phi_stmt_2997_ack_0 : boolean;
  signal RPIPE_timer_req_3004_inst_ack_0 : boolean;
  signal do_while_stmt_2995_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_7671_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_7671_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_7671_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_7671_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_7671: Block -- control-path 
    signal timerDaemon_CP_7671_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_7671_elements(0) <= timerDaemon_CP_7671_start;
    timerDaemon_CP_7671_symbol <= timerDaemon_CP_7671_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2994/$entry
      -- CP-element group 0: 	 branch_block_stmt_2994/branch_block_stmt_2994__entry__
      -- CP-element group 0: 	 branch_block_stmt_2994/do_while_stmt_2995__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_2994/do_while_stmt_2995__exit__
      -- CP-element group 1: 	 branch_block_stmt_2994/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2994/branch_block_stmt_2994__exit__
      -- 
    timerDaemon_CP_7671_elements(1) <= timerDaemon_CP_7671_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995__entry__
      -- CP-element group 2: 	 branch_block_stmt_2994/do_while_stmt_2995/$entry
      -- 
    timerDaemon_CP_7671_elements(2) <= timerDaemon_CP_7671_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995__exit__
      -- 
    -- Element group timerDaemon_CP_7671_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_back
      -- 
    -- Element group timerDaemon_CP_7671_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_2994/do_while_stmt_2995/condition_done
      -- 
    timerDaemon_CP_7671_elements(5) <= timerDaemon_CP_7671_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_body_done
      -- 
    timerDaemon_CP_7671_elements(6) <= timerDaemon_CP_7671_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_7671_elements(7) <= timerDaemon_CP_7671_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_7671_elements(8) <= timerDaemon_CP_7671_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_3002_sample_start_
      -- 
    -- Element group timerDaemon_CP_7671_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/condition_evaluated
      -- 
    condition_evaluated_7695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_7695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(10), ack => do_while_stmt_2995_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(40) & timerDaemon_CP_7671_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(9) & timerDaemon_CP_7671_elements(15) & timerDaemon_CP_7671_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_3002_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(17) & timerDaemon_CP_7671_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(32) & timerDaemon_CP_7671_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(18) & timerDaemon_CP_7671_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(9) & timerDaemon_CP_7671_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(9) & timerDaemon_CP_7671_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_7671_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_7671_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_loopback_trigger
      -- 
    timerDaemon_CP_7671_elements(19) <= timerDaemon_CP_7671_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_loopback_sample_req_ps
      -- 
    phi_stmt_2997_loopback_sample_req_7710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2997_loopback_sample_req_7710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(20), ack => phi_stmt_2997_req_1); -- 
    -- Element group timerDaemon_CP_7671_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_entry_trigger
      -- 
    timerDaemon_CP_7671_elements(21) <= timerDaemon_CP_7671_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_entry_sample_req_ps
      -- 
    phi_stmt_2997_entry_sample_req_7713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2997_entry_sample_req_7713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(22), ack => phi_stmt_2997_req_0); -- 
    -- Element group timerDaemon_CP_7671_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_2997_phi_mux_ack_ps
      -- 
    phi_stmt_2997_phi_mux_ack_7716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2997_ack_0, ack => timerDaemon_CP_7671_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_sample_start_
      -- 
    -- Element group timerDaemon_CP_7671_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_update_start_
      -- 
    -- Element group timerDaemon_CP_7671_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_update_completed__ps
      -- 
    timerDaemon_CP_7671_elements(26) <= timerDaemon_CP_7671_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/type_cast_3000_update_completed_
      -- 
    -- Element group timerDaemon_CP_7671_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_7671_elements(25), ack => timerDaemon_CP_7671_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_sample_start__ps
      -- 
    req_7737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(28), ack => nCOUNTER_3010_3001_buf_req_0); -- 
    -- Element group timerDaemon_CP_7671_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Update/req
      -- CP-element group 29: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_update_start_
      -- 
    req_7742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(29), ack => nCOUNTER_3010_3001_buf_req_1); -- 
    -- Element group timerDaemon_CP_7671_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_sample_completed__ps
      -- 
    ack_7738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3010_3001_buf_ack_0, ack => timerDaemon_CP_7671_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/R_nCOUNTER_3001_Update/$exit
      -- 
    ack_7743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3010_3001_buf_ack_1, ack => timerDaemon_CP_7671_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_3002_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(9) & timerDaemon_CP_7671_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Sample/$entry
      -- 
    rr_7756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(33), ack => RPIPE_timer_req_3004_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(11) & timerDaemon_CP_7671_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Update/$entry
      -- 
    cr_7761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(34), ack => RPIPE_timer_req_3004_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(13) & timerDaemon_CP_7671_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Sample/ra
      -- 
    ra_7757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3004_inst_ack_0, ack => timerDaemon_CP_7671_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/phi_stmt_3002_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/RPIPE_timer_req_3004_Update/$exit
      -- 
    ca_7762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3004_inst_ack_1, ack => timerDaemon_CP_7671_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Sample/$entry
      -- 
    req_7770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(37), ack => WPIPE_timer_resp_3012_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(18) & timerDaemon_CP_7671_elements(36) & timerDaemon_CP_7671_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Update/req
      -- CP-element group 38: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Sample/$exit
      -- 
    ack_7771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3012_inst_ack_0, ack => timerDaemon_CP_7671_elements(38)); -- 
    req_7775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_7671_elements(38), ack => WPIPE_timer_resp_3012_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/WPIPE_timer_resp_3012_update_completed_
      -- 
    ack_7776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3012_inst_ack_1, ack => timerDaemon_CP_7671_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_7671_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_7671_elements(9), ack => timerDaemon_CP_7671_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2994/do_while_stmt_2995/do_while_stmt_2995_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_7671_elements(39) & timerDaemon_CP_7671_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_7671_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_exit/ack
      -- 
    ack_7781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2995_branch_ack_0, ack => timerDaemon_CP_7671_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_2994/do_while_stmt_2995/loop_taken/ack
      -- 
    ack_7785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2995_branch_ack_1, ack => timerDaemon_CP_7671_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2994/do_while_stmt_2995/$exit
      -- 
    timerDaemon_CP_7671_elements(44) <= timerDaemon_CP_7671_elements(3);
    timerDaemon_do_while_stmt_2995_terminator_7786: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2995_terminator_7786", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_7671_elements(6),loop_continue => timerDaemon_CP_7671_elements(43),loop_terminate => timerDaemon_CP_7671_elements(42),loop_back => timerDaemon_CP_7671_elements(4),loop_exit => timerDaemon_CP_7671_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2997_phi_seq_7744_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_7671_elements(21);
      timerDaemon_CP_7671_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_7671_elements(24);
      timerDaemon_CP_7671_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_7671_elements(26);
      timerDaemon_CP_7671_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_7671_elements(19);
      timerDaemon_CP_7671_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_7671_elements(30);
      timerDaemon_CP_7671_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_7671_elements(31);
      timerDaemon_CP_7671_elements(20) <= phi_mux_reqs(1);
      phi_stmt_2997_phi_seq_7744 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2997_phi_seq_7744") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_7671_elements(11), 
          phi_sample_ack => timerDaemon_CP_7671_elements(17), 
          phi_update_req => timerDaemon_CP_7671_elements(13), 
          phi_update_ack => timerDaemon_CP_7671_elements(18), 
          phi_mux_ack => timerDaemon_CP_7671_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_7696_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_7671_elements(7);
        preds(1)  <= timerDaemon_CP_7671_elements(8);
        entry_tmerge_7696 : transition_merge -- 
          generic map(name => " entry_tmerge_7696")
          port map (preds => preds, symbol_out => timerDaemon_CP_7671_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_2997 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_3004_wire : std_logic_vector(0 downto 0);
    signal konst_3008_wire_constant : std_logic_vector(63 downto 0);
    signal konst_3016_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_3010 : std_logic_vector(63 downto 0);
    signal nCOUNTER_3010_3001_buffered : std_logic_vector(63 downto 0);
    signal req_3002 : std_logic_vector(0 downto 0);
    signal type_cast_3000_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_3008_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_3016_wire_constant <= "1";
    type_cast_3000_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2997: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3000_wire_constant & nCOUNTER_3010_3001_buffered;
      req <= phi_stmt_2997_req_0 & phi_stmt_2997_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2997",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2997_ack_0,
          idata => idata,
          odata => COUNTER_2997,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2997
    nCOUNTER_3010_3001_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_3010_3001_buf_req_0;
      nCOUNTER_3010_3001_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_3010_3001_buf_req_1;
      nCOUNTER_3010_3001_buf_ack_1<= rack(0);
      nCOUNTER_3010_3001_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_3010_3001_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_3010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_3010_3001_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_3002
    process(RPIPE_timer_req_3004_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_3004_wire(0 downto 0);
      req_3002 <= tmp_var; -- 
    end process;
    do_while_stmt_2995_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_3016_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2995_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2995_branch_req_0,
          ack0 => do_while_stmt_2995_branch_ack_0,
          ack1 => do_while_stmt_2995_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_3009_inst
    process(COUNTER_2997) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_2997, konst_3008_wire_constant, tmp_var);
      nCOUNTER_3010 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_3004_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_3004_inst_req_0;
      RPIPE_timer_req_3004_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_3004_inst_req_1;
      RPIPE_timer_req_3004_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_3004_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_3012_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_3012_inst_req_0;
      WPIPE_timer_resp_3012_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_3012_inst_req_1;
      WPIPE_timer_resp_3012_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_3002(0);
      data_in <= COUNTER_2997;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(10 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(69 downto 56),
      memory_space_2_sr_data => memory_space_2_sr_data(319 downto 256),
      memory_space_2_sr_tag => memory_space_2_sr_tag(94 downto 76),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(55 downto 42),
      memory_space_0_lr_tag => memory_space_0_lr_tag(75 downto 57),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(255 downto 192),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 3),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 3),
      memory_space_2_sr_addr => memory_space_2_sr_addr(55 downto 42),
      memory_space_2_sr_data => memory_space_2_sr_data(255 downto 192),
      memory_space_2_sr_tag => memory_space_2_sr_tag(75 downto 57),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 3),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 3),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(41 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(56 downto 38),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(191 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(2 downto 2),
      memory_space_2_sr_ack => memory_space_2_sr_ack(2 downto 2),
      memory_space_2_sr_addr => memory_space_2_sr_addr(41 downto 28),
      memory_space_2_sr_data => memory_space_2_sr_data(191 downto 128),
      memory_space_2_sr_tag => memory_space_2_sr_tag(56 downto 38),
      memory_space_2_sc_req => memory_space_2_sc_req(2 downto 2),
      memory_space_2_sc_ack => memory_space_2_sc_ack(2 downto 2),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 1),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(27 downto 14),
      memory_space_2_sr_data => memory_space_2_sr_data(127 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(37 downto 19),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
